PK   N�Xf_��|  �h     cirkitFile.json�\[s۸�+�������v��63�e����р�+�*E��L�{(Y�mQf| ����8 �9�L�K����M�g|���:9gj�\��}���t�,�z�5���]\'�_�{�}^xR47���u7��1)�4�y�)� �yF�vN�LdiV�hr~q5}�8És����K���8q�78�	,쐸cH�1$�z�=�C����f:��ڜ�ϜH�sbL��/�-��ej8�=�t�1-1�9��m���H�s$�9��z�D=G&]�̺�?1��Q�3l~�8��0�G&��icl�C��(���pč��떭ͼi�l5��_	��F�£hQ��(ZT-i-:�EKu���,|Y��8 fq��@���0ۀ�,qjz�%R��b)�A1��b�<�y�8(�qR1���E�GQ<�G�ǗGj,Y>������k,��0��`��eg;�%��_u��#	-^��ED�"�hQQ��Q��(ZL-Y�Eo��8�eq��� ��A0�a�,�Y�8(�rp�8(�qP�㠘�A1��b�<�E�GQ<������рMh�Z�ф�e?�����S�>��U�Sr��4�X�~9[�m��o�:�&��Sc��mA g���S�+0�-s!mFS��aWӧ[V(2:`y��A˅�VQ��5��=�a���.��;I�r��̿ۘ�IƬ�O�S�g K3��4%FH�ei��@hO1�1����f��;��P2��NK�
!Yi�/���z��A����S"K��QJX�57�(˃]�T�<�Dk��T�X�s�S'u�r�EYD�H�[�u8;�R�)}��:I@��ʲ��,�t������]Qz
I�'�ܣ,"l�4f���Ԍ�#��G=��Q�����A��φL�c��(���#9�) >��@�\]�R���4��������w��W�8�$U?��s0v�H��;���?���K�N�c)5r��O�#���E�E�P�u�9���<G�sԁ�y�@�>x +��%�������z��<GY��lu�Dl��� [+��J&<9�VN�ᆣ3���|�L�v �xqd";����h���ϲ%����c`h�HNy:F�Btb�#�ぉ���Y�H>q�����{0�|�q��;+9��=�:�<)B{�=4E;�=4}��Y����O���mݪ��7wo�7e�l��^U{��y�7F�#�R^"�R>E�k��A�gX���E �B�a1Ȱ dX2,������k�X��)��>��Q��)�8�X�r,N9��S��)�&L�͘�Dq�����c�	���P�K5�o��iF�U��:D�N��\�S��@ǀ$<�#"����g��>TY�B�N Y�1�d�+}Y��Bo��п?���y��� ��D�З�<H� ��"H�pGYRJ��Rd��)�RIL.,a��"�r�S�~Xge.yY������))
)LI��Y��9fb�OIx��j=ϵ��4�֪ ��'�-Ca�z�����X��������=����&a���_b�v>�孷.o�P�Uu���ղ[/���˟mg��K���m��*���͢?�P��k��=�Sۛ�>\�&�|��\K�WuF�my�||S� ��yi�K����ZV��o�Z��U�z��v�aP7�^���V�o�9��mϓu����I�fYu�S/�4=�j*$?S���t_�D�˕��h�(ђ�R��`����!������Q��2Ug�b�hT��&M[��v1Y-��-�~����gj*���>M��w�מ��5ݵk��.���^���=��1l�n�^��kW�v�	��SzF�M�EJ��%>,%��԰T:,e���A)��4��g��T^2�R٠�z�_��RrXJH�yǅU�O�f�|;�r���er~�,�]q}�L/���-iƄ6� ���HW(��T��ڜT��}�i1o �����\�Z*���	�"�|��!�-2Rd��K��!������Q��^�D��7����H/	u��J1�I��{Y/Vݞ����sFD� ni.�e��s+�-��r=�����>�xsry��v#yq]�ݞfQX�ɢ �f����riA
k$ef��T��m�to���������q�R@n�h���r+-0	�iy1o���7�,x�5�r�4%"��h*rj2�6���������V�ms��Sؙ����^/׺��~h�Wu��w|}���+o���ѹ�/��k_�l*!O��� �Y�Q�X�)��ψ;@�8�!k�2e�3B�!�iQ�NkAT
3(��0,Gl|Y��!�1e�b�''��$W����a��5(fhV�
7�"0A�A��.h�e渲JX�~{�|h*7Y�n���_&_./���&`n�Y��+��{r�[?�tͤ]Փ��s������MsXύ��jZ���n�y_���w~�L���)�&������>ؖ�Qw���w�߫�]�rU��hv&�$����p���q��ߘ����ɫ�h��������dGA��E3�m�}�3�mښ�k����(��kJ�y�xq�7�V�oUw�vk{3�In��߷ͪv/n�qj���>�9�=��Ȁw�o��;�CFn{mͰ����}wu������|W��Ժ��U���5�������x̽�U�I�`�f��ׁ�RhIO!�q��>W�������r�E�i�Z)t�i9���*N���{�j9q5�D����tvƤR@k9T<ZM!H�L����i&u��$FG�&F�OAzTq5Bz����ٴ��Щ�so!�Т �+%%���Z`(i���E1j�ιF�Ҫ/y�WװP�B�#���@7���̐�ׇ��������F��#5Rw{l���RH}�Ho	a��=�a��!!ņ�%��s��m��>�]���u蘊��{���*缶�������w��_+���!�p��%P]�'=��<ɮ痀��l�a�O>�\��;�j�9e��������ѽES��d��^��$�(�)߆��}wZ�/��X÷�]���C��:�+�?u���2����qF�p��M��]���f""�Ld���03O��.g���^�x/�-��a`�S�o�5��l���M�
J�J���� �q�l��󟚛���	�!W����7��?�e�V���|�PK   �M�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   N�X���a� �] /   images/43b8fa2f-aa16-4fa0-a6a4-ecf006c83c4c.png��wTS�?�FA� v�c ��Hh����*� �J��[E��(V��b���"j�FQ0� ���tAj�P��9_H��1�����C�`8�����3�Z{흇��wn?���_:o��(�@v�n�߄j�P�q{�������������/D��oS����K!����n�hO{������ek�n/�扌���@�B�����0�5ho3<=B��n����t@�a����9*������*����&Ooh����p�8���x\4t�R�`Y�p�B[_T�w�o���,x���M6E���r&�ÅA�XzлwI^g[,晁̈���n���_�k����ZɆ�&�i�J�)�aF^��
��w׽͐�j�-1SwS5fp!���,Sw�<�x�m�S?��mO��
�.|��Tc̑��Q�a�P?����-l2?:�����:	���s��� Z�E�����pu�|5����h@���}h��|�/9�Ø�'�<Řj���/O!ݙ\�{<$�A#��Ũ�!��@��H	�����դb��}���f�:?�q֩ez֬
�UD��'�.�<�-+Vg"�w�v�=<d���Q/6r��<�z[x�zE�]s�=Z�.6e�7�G�#�K��R�1;{�芜��J��њ���SU�@���8�>��R)��]����ak�)_�C��8H��-�k��yBE�^[�T�t<��L.S_JUlWU��`~�����K�.D��h;��+�n�a��Zk�J��Q��͛�ݲ]K|Y���`N��f�6����0<6�vC�c�\�M*T���m|cu�0A���9�$��D�Myׂ,�"Q��R76!��C�x<91�>5w�ƛ��T�SlR���+�f�5�ã��Qw$�j�]����:�0X��f��\���i�s��s�l�7�+9)C5��^��T~������<�:���E�"������Z����Rsؚ��W��ƒ�F��Y��f��ar��I�N�ٔy[&g�2�X�VZ�HH
e��zfDN,�q����3������9��>A�\�:�^m�K��W��r+�11)���nn��k'���"�`&*휶K/�ƑPI}m;&��M���U��i�gԸ.�메;(�Djg
B��	�:f���cT�HX��ѣf�\ʰ7?4���Jb1��_�c��w�M���R����+O�%V���L\9b�x�g�_������d���S�^_
�݁�d�vq�l*�PҌM�+�.�C�Zꈝ�F��9øcN�;"_��aS�K/g^�P�x�!��Aؐ�м�R�V�?y[�C��"��';�I_橏��:U,��F��^��� >�3��9\�y�����������^��2v!b%K;w�3���i�9r�ʂ�
_J<f�N���/�Wmi]��R�W6}�0�ͯ��#�5='�	5�c'��p�H+UP�Mֳr�
��DI�_"��ܩ��.h*Rc�D�&z"�~(�p��I*��N�>�讁�"�܌Ι yW^uV��7/=
c~ڕ�_��&����W�2�1��U1��(��n���j���� 9b���wX�^^�de���&�f��M�����W$4��k�����s&�r�J�ǊD�_��*Bvdb��,2�E�O���ݐ�+�Y�=Y��#��l"���}5�%�Q�=�ߏm��e�\Ω�B7�3�'�F_��gs\ɲv\YC,`�*3����hhg�}��z�y�2���v��_�}�6�L��!ˣ�g8�D��.�5�+l�s�#�D�q�_}r_��l�H(�T����F&�Mrҹ�&���H9��$q8�dlkZ���/�K�VOwG�@�O
S�C�΢�Lj��@�����;�7��034�t�A��7�8.į_:�O$��Q8� ��|_�e�I���5�Ώ�i���3�fʁ_f�)(�����m&���F��'���|Fw��9�m��v��PN�~ r�Ra��a�sVr�Y�B�7������L�D,+�kO�I�ƴvc<0��S��D���K��p,Ah�
�C;x���P�kcQ�O�a靲p��!���x���ѱ#�[�VM�/5�3��¼���!I9��:W���A�ȵ�RA���%	�����c�;�E�δz1������Lr�"� A9��\W���NR�U��=����}��/7�>?*���$�D�c�2��2'�cЁUۑZ�_I�p�r�5�^e��(��^~��yx��Y�Kx���2t�Ne��q�����O������kOyb���喘V:��3� �<�� ��kH���~��$���%~?qC�:B�i���M����hU/`��9Bm�9�
/H��;6V/U�QS'����<�6���FV|~<��1�L��ᕛ3�,D�
}~J��LMjF�d%k����-p240:ԾiWQx�Jc�8�G�H�m��ڝ���W?VW�#&1��'F�5Rnl0���4#]�\<���9?nI{s!�ߢ<<�Q�J���\p3��(l�\��Q��煋�"OxR�F�uB�����*�I�"���7�&��AlQ�H���p���j�����s����0V:���y�m���tA�I�s��*�ɔ?u�#��w�y�%kh�?e����=�C��O��f����0�g�`�����-p��i'��*"Q�`���F���%����JV.§��u���x��k�I���U� 6]E���ڼ��K��S����ȹ�B!v9Y$�n��{�G�Y�+V멷+7�|�C��O&�kb��ڲ��q���у7dI$�d:�+��?�ܜ��h���ŘYFj�I|8*��ӢK��8��3������x��z����)I�����}As%R�1�����z^����X�y���	ϣ�I��n �I��Y#<m��*�_��,�H$�e� �ӆ|�u�X��S�JVn�`�Y��CE#?38
J�^�<������ޞ>�D�U�a���:�IΧ���T��XK4��NI��ɍssδ�>�lY���S�-�*�������~��I���̜����/aS���d��#�5V���A�9���|}z3�k2���_�-�M�,�x��&΅���MkEۭ�n�k�#���N�wcϱ�|�\��>���JE�͎>ߗel\'����.E��ީ��/2�"IJ&�6��{���s�Df.�v�|��o7`#���TJ_̦�4��Q�mb@iO�W��dTf��O�j45&%�2����������K���]�!j��TWǌ���WM0�nx���D��M'�
V^x� {����;��!�*�S &WA�1��Y����`�C2Izf֋�M�z�ą��V ��,n�?�2ޭʘZD����mt,!��ꤸ�B�V���a;��
it�*���=��(�@:k�Q��M)�!=����@�(�r�{1$�2��i�_���LNr�1%M
��`|�j���R�3�b!h��j7��^h�^v��d�[Kd��m�Ћʽ�,�R(k� ������4b[M��wJP[u��k�uV���N��+�I�l��[�!/�T�Ҍ�I9��C?�h�<i��f�$9?�&䈪��aϋ:A%��֪	]�<��+���%&�WAT���i�+G��$"����Ȃ2���V�����z31Pf;��hbC��$�DP���y.!6?	�g� ���J�+�+��6~�w8Pۨ�,mû��8c���W��Z7�:�$��ӇZ�x��\p�~Fj���ڒ��ψY��?��cEs�X�l�2Y�膵c7|k��;���2�K������.��'5�9v�xe�.�4�]˵�1�a�@9-�OW�+�w.Ǧ����SS�4��1C!�kr��$��PQnTOtk���j0"�ȸ���52���,��I�c�Ý��D�#�1�]b�ck��/Q�D�
�_q�s�|���Y`�a��6�bl��v�jP���v"�e$���a�>���7�31�߸��eW܀���n�#��
�a�_y��D0��&�d���b��Q�'���1��d�F��Y�@��e&���aϖô���2�։��z�55�$P)X�{�u����4�aY��n��	�|���	�b���&Y����F�Q]�$�U��cH�߱��>W�W9�u��qn��PMy��LۿN�OCj�&�SW�t�/����EB%�]-ƀ��ߧ#[y�J>�;T)��D&;xqL�����+�"_�w��Q'G�_]�#>�WA(�]<���m�I�u#Q	��oECֽ��<&�i�8�Bв��փ3�Ա��KE���B/������JJz�s�`k�Aϰ��s�>�)Q���h^��1�
�+�E��ɬG�K��=u�_ΊI�8Ҷ��p���v�^�o;�3<�á���uTN�s�k�ql��]�~��<��߼k���y2}^p���W�*�O��`7"*��ޗuun��Z2�N���W(��H��Y�t�Y�9�}#���������@��r���D|�@u9_f�l��b�H�U��n�E-]C8a�?��*�`�q�t׆GeG�+J�aė�1LS^��,E���ji��	�vL��G��F�e!�v��0� ��y�l��5S��0�9#+���b�B��
��@mL,��v�C���yu�Y]�G��I���O��/ƕ��,��h{Gu�=��L��H�cAK�t�Ѫ4v�2���N��f��@7�@�"�A B���g����]f�����(~��^�n7d�"�A.=	\O����,}I�rŨ�ဈ�J+UT
2��R��#7���z��wn�A]��Ly�09� G?K�`�>�z�,�"�L���A���@p ��83+����|�P1'���~p�+�s�	�(9����큒��+���Ѧ���~j�Z�G��x 6�$X����t����k7h[Mg��::S_���6gA�7�j�� ��CB�������n6��[{�#�f&D�sSFcz��x�WؽH�3��X������V5�v�(�Û��IӚάˎ=_��eI=@Og���>\:���H�3�S��c�����)���S�����=iF�o��<w ԐZ^E�շ�r?�)A'�3/��rN�4�m��N�ж�oNI�߃ M儊�(#7��o⎬Yc����BRu�=k�%��uR$���W+�-6t<΁\���2)���s�n��Q�@�-x��h8Gm>�.fٙ-����z���#T�}�k�3o&�1�k���h��������dK'�%�e��ZF��-�c�ƺ�-��З���dg�kyw�53���7 �e�֋9�y�$��ˎ-��ɬ�@m��W��p�7O!���i�W9��xmv˥Jm�=���P�����8s/{�����q�$��x��1�qxT 6m+�sT��Fk�%#��N�l
v K��Ki$�-L@f/pC�:��ƒCQ���b�Q�}nN�Mj�R���C��\��i��ZR�L�el�/�>'ͨ�z�4���΁��!�r�_��n�_AG�Q$��%�Pu߅����L��Xԣ�O{.���cs�&�� 7s�1(��i	`v�Kr^g�E��/�ܑu
�C�����X��N�x�P����W+1�o���E�}�0��?����:�W0�llɪ��so��9󈅭x2�\��'.TUu�#�B?�Vk	�'�b�ō�G�--Q���ǣ�rP<�`�xLk�1��r�(�K�q3���&��7��]�d��kVWM) [���
�ā��Ux�ī�wc�Cp�#HT�G�5�1⁓z�X��(��y���f$�µ���Lz�#~��QMM�>�7����ķ.a�A��T?�53��5'�6d��s�.ܢ��T�F��i;�G"��
:I����t�ؐ}�� Dd�V�P%v��F����R��w�i��ENu/-Aך`wW�~�V?LOC�@f'��VWJ�c�Pص�=By�G��sG�������e�P���0oB/l��Q�]��;P|���yᐃ_R�LҮ2����ծ�X˕Is�n@�M�e'I��ͷ�AlUw��Q��d��"d+��O	`��K�n�R�c?B<R�e]-6Ig�<\�b$w����>�ҵ~��f=V|5fs�G|�-V��љ�0 _���-aCU�2c�Xp$��+W ��6&9�+uz��"H�\8m�z��mT���ֱ �`��{�H�L#���w(�/g|
�)&��k�E��Hhp+l�-;�)M���Wz�&��0�N��I��}��,��"�i�p�u1��D�D3Cn$��8�B>}�쾿��t�W�]�O�<�ߖ��n[�݉ߋU���\s����m�AQ`�o�);��_/�Kc��Jlܬ}����}Jsug.���]��ų�,��
� L���J��te{���0�Q�f��)��E`߻�̬w�U��]�2Au�o4 ��q��:�@���3��<d�U#2�.PJC�|�~�2��L���G���p�m}��'�R�G~��Ű�>SC����<C�"l{��\�H���>�g����C�z��%^"
�t.}��M�����������7(��ɱ��)�sHX2W�٬�����RZ�17^�������Ёi$��ޞ���
b����n�s٤��|�B`-�5$:r�V1P�m)�����9����&����9km��c��{���x����&�=�#}t�?\��<~�YI�^��q,�Wy�V£A�X��a!b�
?�MɦA�7ம���Ee֢��%��'��d�7ېYv+��,���F���Aڱ6�Zo�V4��>zƤx��k������U����[�X@��K��{��F�f��.��HU������2��˒�w06��t"�X���%+*��y��!�Ș\ۺXX��Ɋ$w��<䰖��@��������yG�Z�Cb���2r�Q<�Y�ʑ�/]�
�2�~=��2�fơ�sm*���&���6X�g�~���SN���k�v�!F}}�M���
�S�<�\�?M�,�:R@n����5�n�|H:��Tq�[�hj���s�I����L�Ɨ5�`��C�L�d֊��e�Q&��G������2��1xE���#�#��\�t-j�PW�b|8�@�t*=wE��'�p��63�l>���8��D�>*���<�o-Z/�ݸ�$b��DH@��{'�0�,A�E��H�� ����58$�P�F>���:$Ћ���C*�����\%j�Qg^�u�j���X�1��� ě��Y���.�ڸ����C���N�����$m�P� �x���јFv�{�Vo���2�~*Xg���P�ѓC�͛�Y��v+0`�׳�E��[['� ���-�7�&��0e}�(�� ��c���� �����b� ��d�T���T	4�e�8畋;��A���U���f��=�~�[�gF^=���|إH�F3u}!��� H��).Bm�QEl�x�%4��Qsx����Ee1 ��`��T�g���N�p�������x�7aP��[&����X1z~��n\�)�־yX���Ӯ_�T�0�/}<l�DPȷk9�@�"��c��8u?���b���u��G�J6�n��a��\%�Y�3�q𼤟Yy��Ķ����|�uUڍ�+$[����Y�{���lC�ъ���`%�Y�᳏ ޓ%e�T�+�F���}���Ό�G@b}��-�L�����
�ؖ���g ��N������5���y��� �=�#���.��*�&��7����=3m�8�`8�1����m���m���YF�~��q�@P�$�����s;��'�����nX�b�ג�K���w `�pX@�<s#	�5�f��/fW����v��klǳ�ѓ�U!y��>_/J����z=��_Q����[MA���22��A���r|����j��~J�nS�����'���q���ì��D\?���%�QAgi$��P\K
���+�A����r,�`�S�V�HVy���~]ay-�.�ҝ�����!ͣ��*�w�6&�ʹOUj6*���\a��zY�\�-~L8Y��P��e�ߋ��l�h����-�G�������O>Wsv�z��my;y��T[��	>j@#�����k�|����xLh��rb�.���$T�Hj?Wت�v4�쐼^�t��<xE^Zi-d��Rp��#��r-�?����N1���� 0���0I�w֛���0tǳ�h"�(�qB��c�>m���x|w�1`�BU�j%�ڴ��i��R�@"���!�m�l������u�i�A����kӸ��I~{6[\�����2k\Qѷ̓�mG`\��'��������x�@���^W5�p�2���_��}?�./�r1��o�����	��8�`)� �1�5{��lJ;����>W�T��b��"Z�$V�]J�j�ҋ���f}��&�VŠ�&���)g��x'�Z'��O���c�~c��Co��������/`�ϼވi�u���+Y�$b��ȘO�:��~A+۸(x4~��sr���7D�۷�;�?)��
�m�ᨶ��p�F�{�Lw~���a)@7��:~˩}W�v�W������G�N'l���}1�8������F�����5L���xw~"�|��ʋ��nl�7Ky��?����j�����zl�3�#c��ɮ��uk[!���J�]�o*RM���8[Y�9W��qu}�]�~~o���,�&j����s%_�i�!w� qmV��]����9F��;Z��r�X�(}�搻��66a�"��h����f��M��!uw��K��Y��Yj����I+� <Z���>��Ũ8��X���#��-L�sd� ����s榭�;�x�?����L0si	?�?���t�<���]It飔M^��EQ0�M���浾�c���W����Hħ�������Q���S�Q�x��t��|�m�?J�8�!�椠���
��u�R��w|�0l�f�Ѭ�Bm ~�m����$ȹ:�v2H^~;[�Hm��;��V�^.�H;P�葏c����s�w\=��A������\ �jo��;�, ]�A��2��d���8-�CBE\=y����ְ"�Yg�YH6��
�5�3�S�j@�}<$R��}�O�w�q{����R�~�w4@�q��;#&�/���(*��Y�v`�=�v�Tԟ,��ڈ#�z�݋ �i�Cf�4�?a�iP�vZw�c�	 �#����T=����zh
j��tݛ�������"�B�UEwޒJ.ǚi���8鮌���L������r�rj�ӭM�
��2����?��m����n�V~WYE4���֪�UD�a}�Kn ��u�r�:�����k/��S�I��b3}o�윲s��� ��y��o�����Y;P<t��3.�+�����?SXZ ��|�؍����rc=����|E֩�=�x ���t>���;��&���NN/ҭ�:��:2v>eʽ��j�^�dw;T%���T;�5֚#�:ch�]�0�1e�u�H��N��bB@�!��4�b�<�8&_ ����h� �um���.VCy�05��N�:�=ML��4k�m~~3��I(�=�� Hj�8�{e/�%`e�6/S��~�2�LC�Ϥ)�r!��5}�0i���A��ea���m���%�Aa�0���#r��7��r)���;�v�k6��&� �7�ԍ��!drA�k�p���b�)e(�x#=��jC��2v;vZ��{=,H�:K�Qv(�Fb�-��^ئ�
X�+�૵X�v'X��T��G�!
����q&�T�j�c*�X�5���#!rqZ���&���b�8�wP�gY��K�JS48�`����[��Z�a .�BH���K3������!������|J5�i�Gֲ8��C�	��V�M�6��Ok�2N�2�Y��+xZ��MZ�zb�W�X��\���tf��av�A��^0�'�����k��Bꜿ��{��.�2��%�ev��-z�|�so�Xм A�������𰳌|Ai����%f���������-���Ogr���K�
N���0V�9fVB�o2�]��.R�d�?P!џM��A8u�:s� �	>/�SNv��Ћ��}m�8��C���ZN�г����N.YÜTv�	_����]��$�A`�i������m��l��ެ \Fk���6R�@�kןב�����9g����>���?���հ���cA>��^�������Y��7PR� ?(��ͪ�8���DlQ+�ğfO��
���^�-e'~����㌼p�?���zJ�I�z�ZdW��]��������yQ��Ϡ�&t��Fg���1�@���2��8�R��P�T��9S��_���5+�����f38Ʊa��jO�~�6,0�M����5,*4�l���?<)94���X�� ���{}S���$2��=��O���rm�T�L���+o��=H(�
ք�����j'�	Dݨ�0��4��p�5�Q[��c����%���%C�!�5���XRن�E�w�S��3���<��]FÔ��{�-M;4����&�4<�� ""ذJ��C ��2����}a�J�$;�bz���a<X���x���%�t=�L�;S�-���~������G�8�7yw�쌷+@�Lq2�;��h,2��o���v�T�s�\�7y��L߆��*U�GM3��Q/
���MN�3��7A-�}y�s�Iz@�$Wmd۸2X�����@G� e�E���^��1T�=�������˅���M�<�c��~�e$a�@^����8b�ж~��(1�M�{����)���y��`�u�h�c�ʹK�}�l*P�M1u�7����kS�D X�)^�2��=.خ�|�q�P(	�cg��$ϫliR/��j«@)�))��*��a���N���Of8:�cϘ�.����9�񋺓e�=g��,k�c0Ǹ/�X7��b���� mIl��̍f!�rm��w�x���嫬���m/��o��+c �3��$?Ff4O��`^)�n_/L'u���3o�{�SP[��b5X)��l��+�kߞȢי= �d��{l���'ӇF�z}]h����~N���f����1�X7������2%	�'΅i(��������p��dW�3��RwV}�DP��%�t���e��2f�@'�)�n�q�<�x\*ץ�œ�j��x�s�T �}?��pk& r���bi� �>��p���4��f黝O�<}h|%D�]�wg�RX;���q���j�u�M�����s�h1���Rdtz�t�A׎�8`<����'��V��@?E�.��P�+�%�S$��BU��OHN��Vz���Ϣ�c1�@���}WO��X������Q:��.�?5�f}Վ3D~�8�UBۙ���q�3m'��L~[x�O�/9�b�O�ZәC����J⼙�-�3n�"�B�`I2�y$�>2-54�P9;�뾼����Q��hG�C)M|Ci�m�MjL�/e�ܿ*����ĄϪ��q�ng�K�ns��ä_���ő�s��!	L}!�E0����<l�ʞ&D�ۥ�R6�y�tX 2EA��t�h���$0K!����|������37��{�,f{)g�F
���AeڿD"�%h}�A>D|{U^���	�[�����������Hh��Ao��
*��#�&[b˨f����Y=�v#������ʠ��C�jX&ca���
���DX��ȣ���^.�Ù.��-�G��
�!c��q�s��c�*g�����y�k Ү�=(�`,�r[�U���j��%���z*�]����8��9��{�K���+
a&�Lj���ڭЋ�ucg�Ԡ*��=��������
	�m�G����FA��n�/��>�Z s��?4=Ͼ�E�P�i��>+�V��-0�ԯ�=ivQ��`5|��]Uݱ�NXE2�[D�!\�]�l66��|t݌���.�"6���g#lH�<�Q�ڪ��x�E1���m����b��F G; ���]\��0��Ɨ�z�Q�1��V��!�~X��/k�>; �-�G�����4Su���F���!�������
��e[��j�L�,��,�h:�b�)݆�$_l�j������Ӊ�-kw��UޠS�Y��B5jb�Iڹ�w�h� �KM�2��x0?m���2I��}�-<�j�x��e̔3��p����C�	p8�|�(Q�
��
�O����-�P��Ue��V,%ziƂ��/.]TF�B�#B��{��&��60���eG���e�3����Y=ڑ�v^�y�p�ߓ��Ԙ�Ս�կ���A9�Y�v��"'5�E�^�S�k[�M��Ӽ���ti/_�u)mPW2�.蛅�_ m*(xRiv��}�{��n�?h�t��խ�.l������+�򀂂&#ts,�i�%�������<f1A��l󑭑�-fǙ�Fu���g�d7���B�!5zW��	 �z�H�g�)��:�$=c2�be�7Oi#��~���v�R9�fB��kxEj{K����]��m�hP�ˉ�K�fl��7��E-�kRa���.j�]��6c2ï;�����q�l�l4�$xb'��<�(�ޕ&B^x��s�$\��>V�Eg�&����3��I#�^��ȼ4.���&����Ӻ�Γ�Im�q/�lY?�Y�p�|C�|V�O/:�{8�qK�N���yS��O���t5�J�h�vߺI�0I�Y;8�����ݐ�W,�l9�"�(�_����9Ί�gV��i�v0)ǲ� 5[����U`�6ȃ.��I�Z<)�k_���L���c�!�75�����~g�Eű�Ú�T�����f"�-@_���y�g��ve�`=��a�$��3
��os����I��ys�`ܟU�D�z����L`�__01��7��y��g{֩x��s<똕TwL��Ϸеc���.�C��0)��3\���zsJ�F��*��>�]��I��q�c!��'h����Hufiāo�K�yz�@ ���=|&�� mH�����Ig��c�.�WCDM_j1�C5�;zi���z��x~%��-�imK_mN^5=rr��B��EӃ����$P��d',��1�$)�"��`Q����d�}�委c}�H��P�s��_V�S��(��{��s1[H��!�ْ�ǅ^z+>?yc>_����L��#6;�]D�)���i�.?��M�=�,\	U��˩@mW�Lٳod����9M9�����TX��eCY����6�g]E�Y�9�]�nbi���+���?�ދ��.���_�	�F.�[�����a<�㙒���Ⱦ^�lx*�ZG��&�V���W� �hdd��͂��<2�I�$'�C��P̈́xF��.ˎ�R�/�� Ƽ�%��5���>�.Fm�*�X�n@`f����IR��1�j����	���o��nO���w�s����#�p�����d��]��vz�L<���%�>a�7&�_I����d=��Z%��0� �<A]�H2Z���TA9��i�g��_ f�c�)I���z�с̃�n��I��3X�p�A�C?��͢��bl�PWc���4���"i��L-T���TH���cʓL��\+(�u���:�$@�{��PՖ�stj}������v��'�JI7O;�;0^��z�	�+P[��E2�~��`�`E%�G�]�]����7�lLG�	�,<�e�6�U+g�n
�&����|]<֥�*�������Su 169�����`4.k�3.��o������]7ӟ^8p���PU�&I	G�(m�g��N��M�[g(о.���{ؠ��x���N��7UDM�j]}_��g���d�E��eו�:ι�4;�o	k}�jI�q-�����U]~`D���D��5G��,�u8�vC'����~t&��/OY���I�5=�5p\��2�(X�'x���~��O);rw �U5�nx*S�ӗm���a�f��:Tg�[6��κn�&Uz57��i���t���.'�t�ԚZx�iqNu��l���'u��+u0 ��	0�G����.�H5#��������p30�(�RN*����9h��E�Lr�ڗX&�;�P�F0�9MK+5�1��A*�S��߶��c��.d�K�_K���vdt���~P�F@_0y���v���
���X;L>�c��&%��q�ʄ�	�M��U�<�a�0G�a�K�D��2U쌕�L(u�!t�l��S-F�����Jg3�j3���3�	7�&�h�l����aN�r���{X��$�\&����!bˈF�~��rb��y����у�'�3Q�Z��}��N5�c���M>�ˬ�@�H�ǩ#嫬կE�H�<��^F��?
� 8<[�
�\S�m�w�e��,� �O�@%w���j8⹵l���h��;���H�ZL�$s͌w�.6қ?���cg$'�r<*�2�&G�+��,,�'wֻޱ1Z�c�)�W值�V���o�VS�5�饅��HV�5G}"�0��б��CѤ7�Y�c䪗�<��V]˯tn�CT7�ޘ?7�5��������Ty1�A:+����	7P�W�PW�-Kd�L���@2E@��(I���!9��<ITl�ӝsv�7h���7�8G}w�~��2|!}��d��vZ4��<��Sk�)A
�9�$�Ѯ���h'#�rEו�=��l�D�I�-��XX��&�9{G!e��7>�t��[�5_6�uD^E5��LmH��_/4�Z�U��5����"1��F�:�ܣ��Ě�#,s4s�$Ӡ���w�vE%�v٨e��t����3�Ip������-�Q���wB�{�'�K ��_�$F��b�
d�5"T��;u�����b��L�P��5z_0��T��DEOa���}Q%E���V�Rkα���pR*Tb������0�5
�>�,>����d\8}H��O%?�/UT�`8��F@�E]$.%g^�)�nK����=]pxb�`�aSy���X��O_t����<*S�ҥ%p����w�e��|��DLܼ䍤�/V7�NA^X����1�9����eL�~��l��#	傩Y������n������������Ҫ���0QX�Q�7t{�Ji���h%��"=q��9��HWZ�����\�K	�����M�}� �/�0�����__R�����S��<u5�g��������c��5MC���~Ft�u��� N������Z�-�� '�Kr���xf����_^���N��r�2d�4{�8�����7��3���7��3���7��3���7��3�?�aU����Y���3���_�' ��UA�������\�M��i����3��m9#�6w5���~xk:�{���mZ�����_�:���Tj���G+i̊����4~(A���m{������'xי���c�m�N�ף���ϴ|BM�q���J�{N���x����B��sts�G���v�9��V�X����t|�dPEie������ ٕ�6�Ʃ.��/R���T���_6�v��϶͜�Q��3�o���_^���o����f���o����f��Z�����-�����\KGB����g��>�*B �Z�s�=Y;�0s�\�n]"d~�Z�LM�!
���sp���B���9yv��%� ������n�L�.�3a��A��f�xJeo�)�0�Fb俉x���ڹe���VE���ܣ�ȯ��H������|�+�|ۨ���3ǧ{�ƿ{�M����4�B��P B�]��~`�����^xy��:ǯ������O�L��j�#9�M��7��sAqS.�}~�ￇU��o�II�p�����G�����\�s��7h=|(�4�/��l?� b�5��x�_��	��"�T3�Vn��bw����Iͽf�����z!��O��N�/\t��x�O1Z��r��=�V ��r"Y��R`���9�H<���Q@�.+Mf�����,[��-� ?CNq�m�[�{�y~��2����L���п:���6�?D�R0&g���w{ (H�&�E��J��e�H��j��Z��Q���#��)&ƿ�sS��SSqK��-1@dw:��G)N[��rRW�3�Vj����ã>ICl~�)"����3��aF���|�Js��`�]�(ч/�	����x��uY4����z��n�+5˥��ݤ�-�I?a8���V�C1��[��)�����z至=ʻ���O+�Y�L���zB��Ӓ�Ik����?RۯkWE�<_Y�B)=\=�$<�n������w��*8�;ikf�2���'D� ҭ�����ә�r@;����+u��ϡ���q��?4`�헭?v0�`�y9T?*ν�j{^vP�M۽G�[����Pm	�V�����J��]���;�Ŷ�����?W�6��[l�g��	3�HZ.�qj�> _�q&����5�E� �+"m�W���i�U��7�-S+�5�NN�>5�x�!
�~l	�v��NTQ�xD�
?��A�Ҿd���:r�� �9�ag���-χQ��7�|�د%��� 9�N�!�m��y��E�_L���F��H�)�뮖v�*����z���-�t�����峇�>�<���������:�GJOuo�UpO9���j�<���[�w�5�)�_ >���u�̈��5�eK�+{敮]��~����ի2i�wo_w����	�}1��jr���~z���399�������X�PQ�c��c��QD�t����?�� �����F>߭�ٲZ�=t�|46�G���e{��9t~�4�T�^}��e�x�b���6�����h���%r.�G�ɸ��>�����y-h�s�b<��4�Ҫ���k���~�=cg������l��[V��ͣ�z�P׮]1�&��L:j53�g|�О=Ǝo_�%C��#���Ll��ONH�z�W\�oo5&�r�~��/;ʲ��{��X�T�8�x���}Zݩhl����=����-������7�mds*~`��y���T�����W���:``����@�T��ᤊ�z K��K]EAC_���umñ=����U�Q��G��z0���%�T��Z�	�O�3���t���ҧ0�2��0�@�	�z��6�6�2����g�]t�բ�������G w��&�P�����e7}��2Ґ�i�s�Y7��+eG�Y�>k�m��i�=\�J%������35��\pke�z�t���?Bs��T}�����t_����|ze-]��);�?I�2z�f^���Dk���^�[L�ٶ�$�s��F�A�Լ��RRF����CU�D�=�W��~�m��su�G_���R7�5��*��-�R-��\�s&��?�
�,;�����G�̥{���%2��f �Ϗ򳚆^���nt�f��Z�#Oލ?�)������?��/k]��K�*;�V���+�N,?�%��-�`�{<R}�jC��/�������D��2P��KA@Z��K��KT$�< � �}��C� uh���u������1w�������3�9���޶�W٨�՝�ت�go#�th4��<�l��^ Y����o�n��.���O7|�;r���)ILҳ�p"_"�ɉ"9���;Ƿ����`�o�ن�����������M��m��i�üʗ^��ϛ�b?y~�ӯ�Aڕ�x|y�S_��L	uY�R��{��mwx;��-8�Ms��dPaӆ�άع���\���up�.ʜ':�#r��E�.�(�b3 ���?�D�m�d�w�<�hIz�V��V� q{�t5�����4���򞦏�.�W��|2��qa��� \�+#=��	7ab� ���	�k�"z��쯻G��h}�Vg?���&y�����`�}���J�Ҿ��ł��,�Pj]�M�0��߄��ܥm����!X��Gi�g54�ק^'�s���aAF�w�eã���𪎕:�˨�Ʒ�di�'�+��ֻH{�ps���|�|r\{��4�$>��
�tn�]�{�Xv��2Ť�G�c�Ey�Rh�I:�ځȃ�0R�"����u>%ې+ԙ*J'�ތj~��/+r�vH�a �pϒy��bu�Z�ݷgD���K/37���/p����7a�m�8s��}�Y�٘1���1���J��'6��z�>�H����",��H��#u$55�?���������El�J[�T���+"�O� T���x�=p�'���*������gmz��+V��A�a��$ۙ��.	^�U��7pM�����ĺ�_�b�0B[^�w��㯷])Zt����ik�;S��]>]t�-'��eZw�Q��|L[�6�P�v�­�@�'~N޾;�JGw����]��yOo�?I¿�������'#�I�]� �	Bq��d�G2T"}��miN)���N���$\�V*�zp�'���W��^�����7�D[/�΢wq����耇�L�.V4h
�S��S���>R�A"�E�~�5��ψ��l���	��%�a,�b�]�����`1��@�ˊ����\?jbJ����裠?�Ȓ��j#�V��O�2io���y<a~i�U��rv&�
MO��*��+�v���u���*!�]��+��֘u~�IgŖ 'u+;=w���o���8~{E��>��-�O͖H[����2 �{��+��L��n�Ǻ��U-TU�w.�w;j��8��þ��0�ĭ������#��v��	5����$�J~�f�b��7�-Ҏ��������4���54&vhI3����cԫ��_�0����K�,xbk*G��O�^��S*�Z��t�.ۜ�_Q��Ý��?��o��j����g?Gm.D�_�<?��$�~����j�s��E���0��.-�ɩ'�̌y��2�D�
��U4k��.��aG��ZFQ�����R������W��{Q�,`	Ro.#�s�2Rl��da�6^.ZU�7��В��" �)���MluL_���fK"��ew�d%W���-�툡Y,�a^���X�SV׺�glϟ�	�2�}��֝�����s�a���we�s�؝���y>`#�-���f��
�v���ޢ�xb���)�pa��2Rr����1��ĳ�x|YQY��ǃ�\�՞
�#���G��l��NF���2�p߂t�6���B$���wT-��Ԥ�����Ѵ�2r;���"?.���Ɍ�b��T�Ѭ���?�����庵��d�T��<��� D���37������ 	�t ��ψy��(����9��C��hu=�o�I�s�x\�}a@�� �6qe���������K���mm��)n,:��)��F3�(M���OG��r_7�`�p�q�I���$G"��$��h�K.Dʹ�{��:e$~)|��%M�[b4$��/_ֻ��?��ES�6,#@/G�$�{⿎g"���o:@�x�M�����{.%	$5��z�^M�g�m:�q�Nxa�,Lݑ)��O�0p�r���h�R0�vʊ��1�u3`{��������0ҩJ<i��O�A��|�se����l3�@���Q6��pW��D-�xA�@TOŃzg��F?μ�(����]����ּ��B��cn�-�eX�){%��2��s��lvV`>�(O��6�콑��T\H-#X�L�t�tê��,!,�,AqSVv���%��N:�~����r"���L��&!�
_-� ��t��p�n��0��Z�H���TU_��F���v��&�){+�߿����~M*��Ɲ�U�9������*��j��S	t��3Kf�4ޫP��88!�4���|�0ĝ=���Q[�,�3c5��ɓ+w՝1���ꭦr���>�_��(�:�.qe*ʈ��������)��"�M�d���e�^��4����.�M,�ϸF�>՗��ʡ����@乓3����)'S � ׿��{���XEf�
�f�yĢ�%�� �ג�Z�"����Y��&`pm2��>��:ܫ�6kV�a%;Oi�l�Q,�Z�S�7D>cbRt�.G�UA��s�=�R����)�(�ϧT���̪_���Yi��(+O�[̴�/;��z��t����l�5�R�-�����9��?�މ0>09����M�:f�6�V���i�"�K���Q�Z��|͐u����n���7y���b;�s5�
��gH��T��6�ځ��\���	��L���\J�t���W�Z��B�����;�(O��R4s̕*	a�M T�t ����ʛV|�$�:�4�x8�d�pbJR�M	�-v����͔�l��`�1�:\X�o��L�_�t/�a�����{�,��4."����:E�h@�t�"��G�`���<���3�+,Ԍ�Ey�_y���y	�4��ED]K�����/+����d&-顉��L����Ϭ9I�����"wW�Wɍ�pl�u
�bd��wf��D�QPbu��JMg#��]�7�|��ȭ�Ti�vW�R�%,]�T!�x��&� �O����f譁㚲�%���")rW�Wl����41ޏԶ��@�y8P`����8J�1��$��`_M�F�#��q$�ǝհQ�o�̀!hn�3��Q\pT4���_��8/C���]3_�!�IO/z��tg]o�"��FV��S��p3���jྋ�$��Mh�a��lb���ȵVs��'��w��ǯ������"��T�ӺJ֕����=��)9�}:�U�	��l"��l�tX�Amo>��|���M�;����%�a�q���V/���j(P�cQ�M��?�Pq�u;��q�#�\�`PK�'[�Q��欂;J����i����6_]Vy�QV��b����aHI����V��6�Ar�w�rYZ-Q �a,?IH�Rw��U�ݟJ9%!F�5�b8�#d쉶��u��F@��>8W�[�CSsIl�r�Λ^h������21qXx* F���F�	��a�o�ŝ����ϫ`'�:�[o���qi]�cpđӶ����M��H��fz�M��M��h�n	� VBΛu�<�^|���h�o����ޙqڣ�p�O�����e%����1#���8�.T�`B�0ȀH=�#v�h!�>ծ�4�i��������T���{�(�&@�f슧7v^����1�(�_�W�����p�����AD#dȱ< ���
E��EG5�H�����*�ןί�F��`���� ��7@E��Ti��F�-�+��B��?�v��J]1�G�SC�,�
E1K By�a�z��sܰ?�]Y�Y���*�}��������5C�ڠFk)g��#mZ��)�7_��Ѕn��Ei-�XԮ�9�3�j��p��a��om����L��o���:���j�W�ta�/�fy�*%�}V��:� ��H�I2�S���n�Y���R��bƏ9u1j�f�RI��j*(h2EKx�f(gDR;�T��j����QC ����(8�v߁�t�L���:�~�u���o&���y��i�xĸ^a�K��� 7$9П5�����iO�)�5�x�'N�����p8�]�¬o��P��(&�TY_��Jj��5�T^�5s��i	�`U�#��yӽ)���@�3:D��E�U�1�c��=��lm�D�KII���q�것k@pv�S��	�&�Ux5�(ل�d��KC������!���� �l��+�$��.u!O���ɇh��� î�e���Qֈ$��8�v�՛Cp��3��O���"�6Pb��%)�q��+�&ۤ�>g3��no-fϿ2���p.0�Ū�~��n������!�7��������B����Eۈ_+��ρբ"����3�!}��o7��{�y:�zq>$^�G�E�[�N�O/WO��=�׃}鮢�������k�5ti�Ǐ��W��N\�s���E�������/j:�u�G/����u�x%fZj�,��Y�|Y_�3��S����g+��o�4X�Zu�&�YA�h�=�H7Fv��&�Q8Rxn8ێ��O�ik�����l�Y�[h�?�p��)Fq��5^��JdI�} �^�⌴,?���em3��p��>O�|��0�T7��T8�Bc��`���K4�XMry�p��z�%1��#���9�cb悧h>��Jt}�F���?�ߍɤZ��^>��aR:,$EL�>��!�B�ɰ�A薦�nVa�V�B�W4z\l���-pzIn_9��x��I���?w�9�v�� �b�b>B�ʡ_�@��i,[Yv��Rs�I:��WZ|�'�F�0 ��M�OU�ޤ�U���f��U֖�|4eLBq�Z�#���VH4�]4���wB�ޮKN��U8�F�En*�	�:��婃P��7�11g��DCC���uPy�����K�Q�Pj�2��2p0��#I�����2	���,4)l�o�M{��+	\�G�C�3.n�[���k���ŕ��2~}�K��N+O;]\���L�"��3~�\P}t?��(U>�B6}�d���	�z�$��솛���뙾��/tYQk�̄�J-��۞�k>z��u��bi�Ⲯ��rv�#��3�%\��jpNT
~u5�9�_80<����鬺J�1��?����rݍ��7�6�I\eK�ʏ�3�ji��K�#����-�^��@ ��¡.s��*�2�����eu�\^��^��dDP��G�T���I�)/e���¬�3�Z�3����741�q�Q1�Q��K���U�6��@��j�\��Z�k�j�������K#�����h��B���p�~5,w`"g��Po$4�R�X�g� <g�ܜ�{-�y_FwX� 渘ICA�{tZ�T잞QT�n�X�%� ����FF���F�X��O�-���K�𐰚T>��B�3W�	7�p�jx�E�wu�����! @��}@���|��������/��|��{xU��3yn� �|4�Z1�&�}�+ /���h<�rչ�+1E�)@�d�Lzd����.����F��$$��[\�|�+W�y�H۟����*M6��U��k4�׌��4�Mbj�#�З��MCS���yk�e�5��%:�_ONL���&7f-��%�6�M����yH�!$���BSS=R6��rO�j�5v;o��ҝe��gB/���x��"X����rǀ��`J����u�ї�̝ww��:d�w{���˾�PqӯW,���h�}��?.�X���O��hO�7�����+�^�+�X#;�������e�2�7�C�1�$��3R*�!���*�K%+��9eDLq�pƳSgܴ�V���>��әP��	1v�:�Fq�v��.R|�x��AN�i�_%p8A������k�>x�.}� '�d^{%���㺋�ܘfu�l���(���{&�]��̋�v�*E?������70Z�	�ߑ8��V=*��LRw��΁t�<=����yz�y*a�� <Y�$�]�`[>�|Z8�i0���8�J]0�k��=�FVQ)A��f�y��(MQz&��:�.������aﴧ=�B�".�`b��B�;��r
���4��)̱������5۪8�N�D�3�5gD�+�ӂ�}Χk����&��b;q�n9<�	�-�����;N�^��,�-�-7@w��˖￳����'up�6���p}�˖��w�Rt�\����q�}�N,9]�۷��tu($;���J	SEQ���A���P�#8ܛ��&���ng��~����uE��>�Į�#�m11i}���^caz�Ǣ�i��5�nw��a�4e���,��NL��'"`G����I�nu�E^���������'݃_8y��ޠ��CS���f~�k��1}I�D.m��p峿�Pm5Z�|JdU^m��ZW���Txn�k���nD4,�@zW�ӏ��
�_D�/��/�"x6TPR{W'9����̯t��~X�v�(�y1E8�d.��ih��K�s�Uoo�31�,lnxZ�Fi�[�6����-���GY�{kz�������s&Hzwë�3����A�(��L�H�₂����_Uv��I�Z��B���s�/�{�r���3���A���+rb!7�����RO���A�ԺW&%��=+~����-X�wEVwP#2��&�C�j����ǳ�J����Geb�q��Yg\�/���"ϟej���Γdb�Ƌ���;��y��p-��e0�NrY��ڍ��έ߱�@���Hl��XD� �s"�J��%�,��|�����>��i��]66k5�	UtA�3�f 0�����fl����v��C��x�my|����Y��D�1q���8��!H��x&�7\�)�_X�~�5�-�KK�xӋ�X�
 ��2~��=�r[�&�WT>��q�ɍ��-B�[�?C�Z��&:;��a`�!`%ι*�鷮���c5O� ��ؖ������e�5��U��M_����B�q|_(ڿG�|tY�v�<�ץU�߱�	��@�i\s���B�0Ƌ��2�"p�S���.:��L��O�<�A��=Į�A+��k���>+�R��[*_(�4���N	�<�P��>�s���Xꀕ�Z]������9� #�x����H�7�|CdfT�{k�Sȳ.)��"�V��EM��7��8~�V�Y���M�.*��Q$3�m�lxQ�79�/ʆ��=��M�Ri��'�ӵZa^L/"@h�����;�_Ir�iYv�$�Ɍ%4�jo܂/����YF�X�(ȬjE:c�cQ����I�c����sʞ�+8ԓAV��A��X2�R�X֐�,\��O�g��"(T�x���G���k��@�>��h2��A���Yt��q1�����	���B(�8%�W}7��{���/nä��LG�k�gbo��RyԵ�;�� )�*��	R��q�5�}i���c�')�fU���g�������#��f\��RM��
�b��"��Jz���� u�4

���ڱ/�����\��@~�_���y��}�Hc�@"�f�a��z����M��/�P2/0'�>V�Adg��t֬9�	�g���}�;V�c��C��Z��Ӣ��+����x(�	���v�(|�N6=%&__��>�Td����mY;*s0O=�"y�paђ�蹞��% �vX�`P܉}�O�l)e�ο������$�y?��P)���k���$xO�@@�l��oa"ļ�Lͬ *lY[��sO�}�����~k�~���ϟRS� xg�}~� . ��
QN�Q��q�׺�I,�F	���n0,�U�S��^r��X�n��>#BHŤiG���ƽ�Ìo��>�G[�ʼ�������]�x�JF��ܯ���Q�!p'���8Yi٤`?>f��p���
�Sx��r���d��Q��;����3]PH^P�f�%)�����@���Z�TQ����0n&�x�G�c�p'�\���K�v7���.���╥����o�� ����I�.�
�vTo9�m���<Y_4�~;�F[?�����!�Z��k�uEv+���l�H���"���[5q�E�;�B	�CJ#V���T2��tH����](Ts�|	�ũ<���Q5盶�$RpFc��v����|�1��7�E�M��W\����?��~�~|����I��~���&;��������\���r>�:0�ܐ){A	�����B�i'�!%���m�J� �e[�K��z�M&F��JNSֹ��?�`�)*�k*'�5g`�w������+$q��l~.p�rc%��T �^!vAX*�x�M�LO �/T�����.%`�A��ߛ��hJ�8� 2�x.��`p��~ZW�'�p!p��F��pݾ���H�؅��8�I�h߯LvV ��EK�q�J�o�6�&��=�/��z`����a��W�63��
���Q���`�[�J{�ga��?Y���l��5>?��<�%H=�+T2�uG�ͺĘ$ �;�~�T\�ť럵4��ܒJ�.[����#h߶�^;���ũ��y^p�s ��3[4:���8����ԯ����77
���#ñ����ji>��g���JG��I��Is�4ޙ�����W�:\CXE���Z�����I6�R�w\)�jۣ�%�����n��j���G�z5�Ъq~n��{r�~`�T��_�z�3Lmr��3�|U�"��|�P��2eR��;�8��9����O�V�$d�2�˜����w�\·p��\�j/�Ių��P1t_�n���r�P0?���Dl�5��$�xx��y��"D��?y9%v/�^u��/�]�ng'��J��Z�V$y?9Iw/�W����?�L���j�k�5n�j��	'(��[�V�L���W8���}-J�JI����EZ�6! X�p��h�J���u����� ,m`��q��qN����4���i��I���[�&�U#T�\��]^���|���i�A�p��x����k��R�ִf�����Q�s�@Kג�y<��~�����ĘX���sa6�V��v�~OG���� K0�X��[��X�v>�# ��6qhS���Y�h���)�N���&�O���ZRp�tIj]7�X,L���Ղ����W�'�Q���덪���+*��RW5	�gX>�C&�<�<e�{&`�r�l�ڗ���p(mRğr�p�C��/,��egpM�ȸմP���u�/H�nI�`rҪi���3���1 d�E�`6����&h�>1��wۏ��<D+�/!4��rd�E>�L�sU�c� zX���u2y�!� �R\��4[��vV[��d�aMCd���Ɨ%O�9V���6����h�Z���) ���4޳�ʻg��t�t��$���4r\*CX�uݾ`�C�%@,5�M�3
2�O�? �K�LB��!*�eH���cc썐�9�J|�EN�Օ����l-vl���c�@�V�����K6�8tYd¢��iZdݏ�u$���W�d�)E�آ, �	Fq٦��-l�NB�k2-EOƪ�9�*��b�B�L����[|����De��	nI?��~��ޅ�_���nK���2o�҃�n\�wxoȇ��,��ؼ��{CE�*+�!,�s��|
�����S���C�e�UΦ�Y,�0�A�I�����%ƛ����5*i�Hl��7GE�x(J����._"S�ݰT!=������ڝL�0�X2)އ��G�Faץ�$�������~�ʎb���|�nᲈ� �e_��lD��n$ީ]���:�9�]�L$^G���l�6npȵ%��'>�M���m��C�d}�x�E������"PָX����h�Rg�Ӫ�r�G�^��� �s��'s�c�WלT��/ݸ���� i���T䱖ʕ���|�	���aϪ}��(�!�;�(I.���*��-����x��$���A�V�{��( ?@ED��0F��`�4����!{��e�(���>W�N3��A�<
�,��c�˟�`��@BF�Mo�,|�����R�+U��κ?tĲ��;����<�Y. �ާ�g�=�߉:yL^�|pF]�=� x��md$C���o߉�������_Q�cV�ƞ�:�$�1��8�P���"�|؍�-�Wy;Er��\����Ξ��T�ƹ����n��.�n��^��"@���0�n�*L�[�J{�Z�=C6�Z7�����+`QB�9U���|u>-ܺ�T@68����G�A�q{g����cE2��ԙ���~|�׆x_ +��C�ԍ/���zs��L�.'	ݳ7W�Xb�2^��A|6��3�͐̉q���$ ����n�ck4`��w�|����7�.��	����w�����2����Y�s���k��Kv�Ĩ�3����s߻�.�ۀ�bm�?�O��q�סHQ�	!@i�["�a��\���x�{�� ���!�T9�͜H�7�	_���Jn�eMԶ\ӑ?�Z��d�)����fXl�(��4:)d�6�f��Y�^�8�Z4zq���o���]���֌�	��8�\T����NI���c�"i'� O�	����8�r�]#��n!�������Q7��0�f�������.����"�Jl�_N���9Y�~��L
����bB���U<���k�<2���$�\���d������c��Dw�]�������R���(�<�s6�/�0�ݦ�H3䇊�3J2�Ǥs>?1�F�Ř0_�3��n_P,�UW�y��S��m�0�w�
Td#A�M�5��A[ύ�8#�=#��tF��.����!�WA��;:�ƘN�����#��[��V<e*~��K�Z��hު-���f��k�~�9������3��|f�E�~������cS�[!0Q�J���(�Ѥ�&�db_8*��]W8�Ì�����?�����w��I D�W��F�oّ�ap�{�}��G�f� �h'�ʻ�$�'`g���j�}�tPp�d��ݢt�����X���b�s*odQ�m�5�����*C�0Hro���k��D���/ ���RnS
�ӱ �h��S�Pq ��=�������ǥÙ�����%� ������EA~Ӎ-��2�+XO�.�޹	�|s�
�#p��#��D�P��mF��a����ͨNv�!.�T�;0�w0��_�'�|`�3���F���ɟ[���܉d�c|'R�ti5Shc�5P�<�3�����lk��h��Z��|���i����}޽@��4;a�W��4�ԏT�upa1h���f'�����웲���q:Ѥ�ܝ��Z��q�
Zs�p��aIԟ�IMN�y&Hu�~P��G-fϏ%w])����I�Av?k�{�ǐl�+ND@.�u��=ax��_?g�,*�k~�v�^�g�*�㍖߈�邧a���������ò���#�ψ�Ty���o���H�A��
6s���먲��~6�ԆWTO�d]Q
_��:��	K�����b!���:a;�ЎO��LNϴq	����O�SN�Hl����`#�^�]������M�$���
��9O�߹+KMP�)ꨢk�q�[��Y+#:cl�_cb����jg��K2�Z<��`r���q��s7���S*a�pl����'��^S��e�C(�3y�����8�ҰtOz���)F�s41���h��j$�fXT1�N�K�|�z'5w�'�H�drR����]�޵�k�b�X'�6 U���L��>1��G�vI+�lQ'�C%'t�*�w���w��P덐Ƣ\(Ti;CC�:�'�(�1?��f�W�A��<?ZO�D?̚U�\.���{T�X������J��Z\l�l���H��N<f���@�ٕ�Sɥ��P�M:�ȏ�p�����C5]<P�v�lv�C�|6��rr��΄R�FE�{����A� �����sD<���YR�TS��Y�O��m]m߫���K{hx/ >���D�,�u �x�[�j�I����$>���xF�y*^D������Q*��F�+BG?ͮv��/�#��Zh��;R�� �[;U5��l�}�xi��T!c��q�wO'(.�N�dCR>�*�G����)��2�c)G�ч$��:�l#�@����!gQn�Uꇮ���)�d�^���n��˰Q�U"ʫK�~|ʛp"oZUM7���;C$%s�5�#���bئ�Py��qm��B}9���%�35R58b'x&�"�_���ʏ?���gg��4���m�y.������p�T���i��>�/�BEc��M^ (�Ff�e�$�+��O��n�{�7����G�l�t�2���x��vɞj����EU�פ�X���n�c��"���f���u�tk� ��q���z��G���}������~�?袌n5�6�GJ�r�O��A=�DW�)ȹx2��`��e:ͽ��RV_t�����|�����4��ѕ7���/�TY��ږ/P%���H�s���3�N_�1����7�^�e��8Q]y?�io��l���L�[�Z�fUyaðqT���g��}���Oo���t|�[n/��)$c#1��K���kA^�࠼�o�~�[!ޥ.s�9\)��|�t�\�%�c �
VK�u�a��ʨ�� S�B���O�P���3LL'��Ԕ���������s\�:_Gb�W�S���j�����mR������-��p���.�-9�ώ��G,Hv@ޡ���M�u}�V� ��\I�������'�q�D��*�|	 Í��`©ca1���A!O���rˮlS��v���~I�*߈:>��OM���5�`�)��ӧ��}�Su6�J��U��'X�\q"�\�':�d�0>Jб�ù���t���PYqX �+_��E]7�(k<�Ll�N�l��cfHW�����?Xٱn�=�'f9yw�ݘYT��c�7h0
�@����}�W���'Α�y��V7ì|�gd/<���-�Qr!I�UY{�.�0�n$�}?cl�Y�V��tϗP�$����X���OϦgZ�X���1]g��ۼ� ����])�N�A���a�����%U�t�fE�K,;���bnu�(� .���8*����t�}v�ۍ��l�i�����+HY�}E2�P���� �����Plt��`^Ue��1�D�צ�2�w�����{or p�X\���c�3�`����>)�p��|��I�c���X>m��>���� ��p1w�����o4�k47���1�n�{E���/���{�l�;pmѻ �@��2��/���˸Ͷ>�	|���G���k��/F��K�Ao�Mn7�>{�[�T����gp6�-bєY���s��4����{T~G��b�5Q24l�����y��n�:^&�TSy���5�]���
�D��3�������~��/�2)w�Īd=:)ɜ<~�r6V��g��[�X�	���F	�f�,CQ�}B�����I:��_�(��GX.,�"� �c�ͮ�K8��-pJB>�*Gu�˂�O�n��+o������Ȗ��D�
'P�J�g��+�l���˜(6)��7|f��.-Jy�f}p׬K���ܰ(�ɛ����\i��ϐ2N	D�[�;���| w��f���ցT&43���3UӚ-��NϳVv���t`�e��r�7�3"�ŵ�߭�q+��r���~{��@���E��ڽ��%y���?�ӳ��b(#,~�_&��>�ɻ�;�$��>j{ȦJ�-C�[[��b���yۢ��"��v��K-P34�������l��(2Az�7@|}J���Q Eq`�Sߐl�a
H?�<�:v��e���٨ݮ|����\������u!t<D�5n����Ξ\\���ύ�h4-;¥o�F�EV��e�S�U P��X.����RlZ[*=�m%0�N�N�J�	]�9f��$#���� ��|�Ah�6o=�?�ύxv��Z(Sa�-����-/VU�d�~�����ɸ�0Y֐8��CU.�ε^��^�:z<����Y9O�e���p��8z]����=®�HffO$H��W	p\%�&�Z���q��e(�<�����2"<:;�ta�+;YkKl���G_�Mǈb3hɽ������'��#%$9�r�F�`���~���4�C䠯��XmD*S|����kկ�v��X,��;Xl���H|�����F���`@ˁ��ӽ��޻��#	%,��t����m�����gu�V��xJ'���]��8�b���;�[&5'�m��g����Dd�����^���h���v���67�y/��]�1�dZ��$0�zn�`#r.쁼�G���/a�

/�4sy������H�.�E�i�Q�N=I�};Ls� =�i!!��w`}�v�"��
�qȁx/��$*�;ů5��UP�Z��J�}��S�׷PK22q�oӀ3'&�2���5�ѷ��2��l�ݵ��h�ί3�5�F��a�}Gס��d���2N��?7U;N	��N��x9Y�g�x<=�]�0�p-���⁖-�JpV�xO	N^?A�:�q���E�m��P~���KV�BP�H�{�������G p����Y5ed��_G�b)۝.4(i����S\}@�4t����H��N��k�sؠ��;&
/Q%���3"?L@l��]���M6�2��&EM��]�>���~˃�Z��yN�+l�|��D�k?-N���j�<~9�E��M�i ��NEr�#l�ߚK�]sӋ��uk�2���|��oo����X`�X�iIS@�Lo��(����-�E��Z�1��3��u�
����ñ�[��Q� f _^�?���⹯�P's�-e=����jJ�ǆ�?�p��<+?w�9D��#!�׍�U��ԟ�A��b��x�|�p|G��[G�N�靇��H���|���-���Z������#�3�ӍM}o��S$��n}|^p��! h[p��k�1;b���u����=0s�7���@���<���j�x�#����8x��I��K���(��@-��>��i��{�bS��(���`Xq�����M\_¨ND��)�O�����_Id*.���b����Ӛ�j��N�}p���?��גu>K? 0����)i!o+�&
����o�	����>Ҳ>1��V�S:f�z�e�|9h�%h���[��eM>�j�Lŉ������I%�� �p���I ��t.��.����*.���ax<�cƱ�tN���$-�ߏ�e��a�Vdqi'Q��u�j��Em��zsi�z>�,�y�}�шKJ��o>����܂.k:��v	���x�@���5������+��:	x
��&	�?)%�o_~�1'�g���qj��aA[ȆZ���c��C<�·j��%�Ó��a ��EF
���2T��� �*�㜥�̛�.)��>k�vߙ��tY2Ay����B�Ӯs��_���N���Ō��@(��vx���Yjk�G&����9u�Mش�o�Ey�!2��� |�7m�_�ǟc�$eCKr�I���ҍOE�n��1��W�MN���rEO2�d��+v�/H�}��u2և�a�]�G�r3Q}���6�B�&�,�'6��
ل,�;Rؔ����O)�>&�Mς��� �z�F\́�Q��Q>b�]�
KpG�W^p��a0�O��4���Zw��+�V�W[j���p��@���Z��,�]���D�Z����T����U�%JFF�L5����E����{�{'و޿qR!��p���_
[SǷ�7�pR�����qF��]�5��)#x*�c?�-�PZ���V;yMfx�^���4���'���\ebX�M�C/��q�ݝT����_-S͞:�&Gpt4#1�ީ���Zgo�'>�~K*6��+����s7�?&��5~���;K�����o��n�@Ҳ��20�(��f$ �+���FZ��{�X���޸+���1)��$z����������{���S��@���=�rtቋ̓ �GU�B��Ųa��5٦�����#�g|���ep�w�;=�|�?'^�G�{�,ۑ�;myܜ8�{���)��p�%[�d@l��ؐ�c�IC`}�LM��Zx��ϙK��7Pa��z�H�󪫢D[����e:L@}?6����&"��j����CO����)��p�yfY�wl��0k簿��#a��rM�̿f1 �G��k�U.D*�<;�!��c{j�-�3T����VqɟÞ��+(�Q�E�Z��`}[�^C���}�X����v.��EͲ���,����f�Q�}Gg�?an2.���D��B^�lP��slx��v=@����`��1ŉ ����g��zG���U���j4�H}~���V'�_@�c��	��H�s�.oN�n��2dײU1k�yA��$A��W������_��8$z߱�����^�x�	��>m��b9��:�,��tF�ߔ�M�۔�tIT��������]��G��>b�G��^nxd���X���F����U�F�EC@%�|�Yn��ƒ��;���� ��G�3;��~[��.7������w��\������ҳX�ۛtQ�閿�x�:{ok/Ū��}�TH���4�~_��ل��r�?g��(}��O�L1�t~i��kb5Z����]g�����*�F25m%5�ͭ-/1}�
 i�A�#�����*j��^�i e��"\t���&V-b��䃦�m��ZؕZ�����؋�q���bp���Q�N�zs�����G�,�|�R�I��`�va�� ;j�W@�kR^�թl�הP�Rh]�^��H���=�r,�謻��3!�-��J�e<4C��`�w�|�*2V�������p����Ҟ{���'�`#�����~gٙ��1R"�:YY�G�2�l:��.���J[����z�"���՛
��i��Mx������=�<���[-WFhC�D���EG�+���<�\��fT����6�$�NO���Z޸)$��`NJ�i�5ϭT2�������}����ȡ(�f�Ȗ�RVn�@x}$D{�Y7$	5�?�̙��rC�o�~:����N�eQ��=4���T�ı=O��>���@�x d/�B��B�g��5-,�Ǽ��g�F��D왳5c�e��͒����6{[B�h��uX] )�6a$�qݒ��g.�V���~�J�uk}��T�6v �zk0wgf�_���f�5�k���1ة��s�4FX[�J�����6η+���J�~w�v��׃�rͱ��4�.Z\�Tv��8�u��
LY�V$��c����$�?�]y��0>�y�o��`�L�̆ä��p����\�|D�Gp-��q�.د[�Y�����R��Ci+�h��9�<K���Rv�����Hm6����d�^)~O�-�T��)�!�Ë�[�ʖ�ݧ����fGR���\.G:��23��A�t謔`e!)��2�#1�çl�����?e��%���ۇ��{���DMd�Bm�m��T�~^[V��Nh��4��o��7��Gh�[��͙�u��Ƭ/�?�[qL�4rH.�82����tg��g��,�1���̟�`�~�y)bb�+v��>얤��W����j[«vݦ���cSR�d�P���F�C���/�䟤�'�o����h�j'�Xz>W��^�z$^�QK��z�M�7��P��۠��jbYv���CG��ؠ����߯x���t9�����Š���������F7 <�{�\S�:�y��lˢ]H����C�/�l���7E�.��KYB�VD.�L��#�6@�� �?�Qlݾ?Wa��U{���R�i�ʅ��N�u�Ʀ$|Ɲ��0��eg9�0��)�j�]��f��~�zN�UQ��!�ha�N�;�"���1\���i/%?�{� ]F�&�KJXI[kz���ht���
G���T��+6���F�1�{�p��*\��'X�ŗ�<7YE�r�?�IU�����+l$6��.'v����&@�1AT�����UN^e�U��?����/n�w���^��ڷ?���8��P�C�ҟ���k�l�b|E�?���HW�"�z�`�mzd����c{ǩ�Gח�C���Ouӭ�����H�5�XۨlE��"Fd�1v�+�RY� B�H����,��%{�:�ƾ��9t}����^��2�s��,���<��+
�R�s3P�%����a|ޗ�5�������E��'2�x֙I<���\�=`Y�lҽ��?`�� �ď�R�"o�C�T���2s���ԩ�{�Y9��d�U'R|B8��;cm� .B�q���|M����{���.^љo^eKỆ�v|O���=Y�n{Cׂ�����B�� e����Gqݸ}פ��_O�
��]�v(/?�gO��J&`�*>Bϐ�F��T�o�3��~���E31gi��O�<l��;���.���m}
�V����u��(���%5�]f�?/� 78O�6i�'�Jc�^�Y ׸�a�q'��n��;�&C_a�9��{��[�8t��]-
�Σ�V�]��� %_��Kd��/<����a�mf��M�q�s8R��b]�:2Q�'��Jj[b��Fiv_�����Kgmt�9&����>��H�:����׏�Z�`�����v��aveh����2�7�X�Q�?E�z�H�Nͳ3�f����	A)ʉ��Y�<���� |բ���1���܈Ѝ�]_�oO�~�kGT����!=m��,nz�b�y-��������"���,�G^}�l��@dǂ	��x(2�5����/�'��=P��<W�� )u@1�����$�Ҟ��fJ!����zɹ���শY����Ţ��7jL30�P�V@�������KE���P�����W��1G�y@�R�\2�l��}���1��H,��X�<Jd�#�]��FXY_�߆p��4����K�6O�su�!�؆��5C����*>�t#��}�����Z��Li,1�4/�W���،��!������*����ZP�rք�o�q��J�������<�u@qJ�doS��b�Kz1�(�������9���L�(�����X�m~�6��t�ϴ@bn������[!���7�z ����4�$�I--����o]ѸbO����}�����E�>�9 ��I���sI�V������n�@;�Uvh"���J�Q5G���fg4W$N���̪q�`�M�7-�/!|Iz�&�w̔���� �ݕ�B�h�s(��t���j�����1�V���W�^��7tγ�����r-M@��]��c{3EK���\��AS���;F|L\�Q�Ŭ�V''�?���wúU�;x[�AC����C��7(����L	ζ���Ϧ��g���F�m���]N��4Y��@C��V�굎c��V�8��U�wP<j�����(��1eឈ�%�El�
�d��W��f/C¦�8�* �FJ�l*i�?e�x��t�P�`�MUh�] �B�Z1=&p��8�:y�ڦ����ʩq��7B}��W�cݦ��|$���x�D��?u~Q�����i7��_}����=������	频6�����K>bb���ʽ`nT��?�*@��3d�lS�X b��<�:@0_��a��T���j?|���WMӂ������1 �lT��a�'@P��jH3��ܪV�&��*��?�����?��	�ץP��c�pԠͣ�l�惢��z ������ީ͝ȓ�RX�@6����?Y���wh �U��ҭ���
����r��Ƶ
�6 ��Q,�L�w]�@�W"«́�q�_R���!�&&�a7uc��4f�,��?��۾sӾ���EE��4��2v��[`��E�\�|~v:nSP!�A�X����/{W�o�Aj�ᠲ��f�U���n�o��n�qvmv����8��si��"O�������or�#P{wI�Q����&#euU���/Eټ����qX܌����-�&&����l�w;>f N��k�Y�r��;��O���?>�~�l����p��߮�`�������,S\�X�Hqs�F�<�/#{7#z�y.H�f~���Ȕ{�¶|1z�ĝ�!�o���0�ߵ� O�Q��������y6=5�����N�]-���Y+���N��͔�:�ɡ��ő�r�Ij{�2u�������P(~�]4�.߬��C�~�	�Eiدh�d�a��S�^�vSsY�d$�������!��Kt ��$�G�l�U~�ґ!fa+$kǬ�r�U�3K�3h��\���YE���%��F�U{������T�yT���uG�c�O867[VE$�<q`V��t�5wh�j{���s�C��V� ��<���5�H�q����=> �F �K0Ӹ(��{Zl��V|�򳚿�ΞKr�H����!�nIͺ�9Q���꺢A�3�.�ioь)9$��u&�K,##u6.DܦH�!2��l����'�,��4p����	Ǹ�k�[u/fZu�X��%ǂ��ך�,����+�Qeu
cK�{�-�|e`�Ň\��&ĻZY	l����rʉL�(��c�3�uѝ���Y�hu�)�O��9����>>����YV���C�o�Yt<Q��{�ۑo�|+�%	�ۈ�e�[k�.��g� VF����ps)X�0��0�!�)Ƨ} ����ɥ����n0<4~_%��Ė�Z���e�I{�@�P=/ʙV4u�`���2D���j�k\O�vr���G�`Μfx��f��1>麄��ba��6���U�^b �s����0�)bJ��0Q�\��fK��[�3l���c�?҅�zU{����N��'ׂ"�Ө��5!�E�w�T���c�P4�j���י��ڙ�v,�$����
d�Ȑ���-7��*X�}���#ISnY;F�t!�:�uX/gj��Y~E�Z�3�@C2�A���I�i�����f�}�@�x�<_�*^���4��]�O�/��;ǵxˉr��A��u+�[z-�i��� ������[�H�rZ誥�勱�Y&��aOm�s��-�*���Nɴ�N1GO>�´��h�]�sD�ݏ�e��$�#_v�O)�9߾x�AD<[��xa�1j_Q)�[C#uG@[���	�J����x}����(�w��t��y����"�n:?L}1��*�/�%_t�*>�������Cl�ۖ��#ᑱyl�vYO��瞸���>�����nT������P~��L���n=6�
�E�Ak%�P]��0,4��>�.��mBw�*�0���An��D�o���Kꉅ�/��n��@!��� �M�������6���P�n����bÒ��+H��k
愖6�@�ﮡ2P��~����E��\L�Z۹#���C�v�5My�_��Z�ly�Fij����~�{�������:)��N����=!���6M��@���{����)���J��h��ZW��YT�@��������=U�%ҫi���#�M�Gv�āS�2�ߥS[�u2f��I��y�#]�{)��c������Vc�LR`�Ò:���ӗ˾� dS�.��;��0���� T�w����r ���󶭗_��\[���7c23��Ҝ�;�L�)�k�f�V��Ut!A��	����d���y��-܀�r#&2`�����(�e��+Q�٪�0�pz����k���������R�o�BvR�-��]#;
b�"H�\zK�>�s5H��hm.t���+�#.����#���&�_�ڹ7� �6���</���a�A�3S�%�����h1�vG������"z���\v���&nQ�$1�O�C�+�{2��^9#��1q-%2D"#�o#x^4m�5��R����\����9��^l���������J�=x��X>��No��wʁn\�Ǚ�٧�d��YGw��i":��+���,QW��`���׵����0j�,27M����2�ب��������� f٣У7��[/��V��j�I���ad���.ZM��E�K� ���7j�C�J^&�ܠ�Uq��>�
�y)�Z¾��5�\]� ��A��;M6��B�zB�#�c��������
��	�W�(�Q�S}��ޅ�u�oS�X=��q��F4 "���֋�Bø���ƺP��`C���ע����S��C���H�� X��0��ר/�x�J �8���Z�J�wi�BWH�ҙ��'�)�-�]r��1�Y,~�.6�j0����	��i�|�v�ׇ�hu�k�`?�j|��)���!'��v�{@���hF_��a��1)V��Ҩ+��R�d�[zn@i E���g@Ͼ���&��]g�EV�O%����b�a��|�/l�|#ׄ?H�$^�q�]�S�n���k)U����ʶD�#�O�}���sڿ8"mQ�U��)����g��9�����ٶz{���|�H8Lp;/��(:�Bj�K�(<d]����<�NՏ�OT���O�9�Z�e���ōQ΃Q@�7�\�b̎�C?7��g_]�+�U>	�x��F(��%�Ʃ21۱ �����(@Oy4�v����.�m��%�n��B��/�- T�ؐ���n�|7V�eu�zl*����-NO�=��V^wA:�a;h���_�5�=�N�у<�t޾��aP��^���qx�"�(���p����;���5����/���LY�e�+�^2��A�v�qF��K/~`֎:4Lb�q��,�>' -fk���ҭ]�F���w��[5&��[+��[�Q�Ɯ�Q�W�>���up��m݂�?�4d��l=W�7�K��K�&�e `�Vф��0o��@o1��P���"D{9ɀ�%��|���/m�|)m�ϠAP`=ߢ�J��'�և�j̤/[[`��=s�E<b�@W=�  �`�O^^�ow�w�匀�a%��%ƿ;{?���}��ftz�}�6�-��_��l�<
��z��H�+����'E���%R>p�+�QLR_@w�{ydZ-[#�ю��1�Id�`�����!�z��:@=�C�Ô��/s��B@�,X��a+?�VcGx,kC tX(B��r��}���<�i����f��5*�����bG��থ�R���%�fn���]�L�y�)@��rO���5"Ѩ�n:y�2sp�a������=�Α#,�^y��o-!2�dx�~Z�b9t�i��	�n��,���QJKu����o��L_q]v��P]��H���\^p]Zj�Yw�>^�%F[�X�hm�jjy�6�2~K。B���?/��t��n>�ˋ�j&��D;�e@�őW���
�nH\�����x�e����E�Y���1Y���E�%�5�jO�*����cQrs�W)���*}��'��a�;1R����0nY������ L�V�C@����m�'�{	�][K��v$��EUS7*m-h�&p?? N��q`�X����r0����)A!��m�g`�D�I��EZLk�_���8�ne��:Z>�1�T�7�6ʁ���D�JO�'[q�����Vsܼm��R"^z+z�����wP���ԯ K��b����@v�(d��.O]���HKe����F:ri�$����gIuN���c	�sȱ.B/G���ֹ�b��E<b�"�y�q�>"�������l�!��0�"z�:*k<�⎵-�!��r��T��86�YA `],���Ԟ�=�krJ�ΓNKCN�O�5���~�(��0��|��?ΘNխ@�����D;�$1�'��(,�������tv �:�����AD2KS��a�o&�m�yAIZʽ����_�X�@���0`=7n��Y!VP�b�t^_b~������]�:���;�j����0��*[{K�\�؂*ɄI��y���Pz[j`&��/ �Z�>Q��:�����Uzi%�,Β�
�Ӛ�0�8�p
F5�ɟ�C������;�[�=���>JS����.�������p):�šxW�%�m�y��5����#�L����8壭Ν��s{!���7����	�'dҎ2S�r��;��8v�N�:�!�S['2q�.Ad�$%P�pat��B��O[��ڠ 	c �;9�' ^�-Yn��X��"�[���|����؆C1��4�ap�Q��c�pG���8�18~��0��k�T�$A����ƩD_�0�}N���QOiJ��aG%*�f25=K�z;�,�{~�O$+=A�-H̍�D�����0ծ�|!|I =>�������*Y>�,�\��*�_���H�� ��S�V@�,t�����G�೐�P(%f�V���&@���?�Af����s��'�-��>��<�����@���筑�TR���%2�7z�kV1�F��`q���U[�]�d���2稧8�����5�x��YbL�9j��:Xw�>���:�gC���;X�bz�Ji,�[/	�j��z�~�mP�{�n>8Ѻ����qs��+m
��cY�������v�o��Rz9����l�pXL�Q��$�Ey'�o�#���6�A��r��K8Pn�=���O	���Rҍ��=G��7�CUr?�}�;��F���"���`mF���Jp�6oI�/��T�Nʅ�;�!�g���l��F� _؇{��������C��q�����/��08]d��d��lx���\�X���^!�	��u)p�ov\&nQ'[��:��ՙ)��ؚ%	� �݃R<��e%˟��DnT�I�9�-E���ǘ���6ڈp��$t� �������,\D���rf��f�c�)u��~����� (l��A!!�U���5�8��]����)+*@4���'���t�,շU���l[���'��RNW������B�����5��
_�����0}�(�N�=-{ �߾�J�e�t���c�ۨ���B"p$�.'GD�#�� ��B�4\F�I�M�������-�Ϧ�x�q.�; ��tނ�q����
��Nd�NR���!M��pC㡛��x�Lh�T�.��g��j�, �åaċ/H.����&�Hq�&�%2��1�(�$�o`i#�ka�/����\n��MeA��}@��ߍB	�IaQ%����Y��$U�xxE4�ӣc�`�#��吖[�Ǝ���w�P�q�-n)Kr@9�@P]{t�ZGƓ+�^N���A�:cj��U�]����9:����8�c
�NC�{�09�v��y,�a�N �6��y���J��k,q`���r����w�̜��� ���V��\��S0��BlC"���ܟiy�0e��j��xO��c忶Nۿ|F
�
X`$�j%�P+��]��� Hh��?��5��t����A�֌:��}�D�S�*ˀF�t���h��w��5i��4*�	�g?�
Ȭ.�����r�HC��T���g�佾m'`
!�
@�q�`��N��F�6��G�I��L^���t��$�GE���9��]���܉Y�à����#���ս!*KHW�>��q��q��s�{B��KɎs))�3-�@��@�]<�Pl��҄^�x� @�{���<xd3r�ۖ���ua���!��Q5b &�(��W�>�{��k�h?�*u���l��( �Q�[�~ƒ&�����X�'���_�)ݥ��z� ����	�,�f��[��=Ǥ�������M?�����>pC�?|�L�JRLJ͑�{3S�Ѣiw��h���ݩ��sL����`e��Q��,tv�m�a�H�#����l����d���~k-�]ܘcdM86U �X�T���3 J�p&�ŭ��⨿�T(+���v:�k����
)�rN�o�+g��\j��>���x�/�A3@��ُ��o�^�� �~УB]��g�y_�`��1�}���kk%ت����s�ioC����� clImk3�!3[ ��v�V�� ����c���e�'u�c2 �e-�"ϼ�yb���a	Y���
4����Y�]�KI"���5S��{�ޞ�Z���M�ɹ4���)�˱�f�Z�499�:�w�6���~7��:�M��
�:P�ڵkN?yǧڎ�5��Q4E��ʐ�
��	����.i���N�?
Z���6�9�mp��qn�����\1����Wf�in��=�ɾ�̙�f���_�>��D� �p���z`���&H=�3^|&�/b߶U(��%/uJ�Vj=��K|t����g����N����5���ь�[ַ&�Bބ�%��HJϸX+�Ho��?%,C��T�v�������li
f֌�:���9�e���u+b�����#�,[������X,W��"�����UI0���<�����񝬎��ʇ7niG�s8,}[��3I�K2�>bu|�������H,bS�����1��N�_�wu6������R1:0�擎���I,6nm�j:@���OWyS�a�/tI-��?���G�����~��b./p��jѢ&g���ڧ���/��G��+��������ic���8��1|��y���|��o�[R%�<r^�����7Is%��QGjR��'/tl���=�
o̩+���"��ߓB2T�r��Xf<���Ыs�,i�hA,�X�$�I��b�F��z�yQ�7Q͚A2���^�n����I �-����>a��y>�"Mܕrs�Z�)�n5?[k�Ou��y���Ē�.�n���_�&0�n��g?oN���Ƥ��s��`�/Rz�PBb�	�֌��QL�����>���k���Ba�s�N~��gK-�Ĭ��: ������ �9���0����$��:�&#����e�G�;�=ײ�q���7�PCz ����>u���LSc��Ϙ��,L���׼�~��i���33Q�Νn.%`.�_S�)Q�/��C	ؘO��
���ts-�����M��S�
�ۧ��Ko�����l��\<\J#��+�tYA�۞�O�����!����� �?X~&M��N�э\�vw�q�8�˷ޛ~�=(�\K7n�7W�/����Y�.����LQ�7�� 
��s	�wY�� ���d�J��s��d����ş��+��j�/��%ej���\[�i�c���΃���	9 ?�JN�<Ȗ5��������/#F����N��Xj�M�B���In�u�<d�L������}W�G�#��r����|�vo��v�����N22v�[�U��ݶ`�ӭ�$�l>)�V�}T��^��2�9�}���7�L�:�G�!��h'
ʍ��+~�����ɦ�X����v5����
�������<�6��8o�Ea���V�@��m��l��S�e���n�s�3({��+*R��ca�u���.]$��E]��{6��Ǘ�Tu�j���Sၲd�`��*v����8(00��Gk����r�7�En��Qх��@t�5e���q�>;ܜ�@	2�x�l�(y���v�C쓹:8��U[�`�z^��	C���m���.�Z��C��l�l»�P���P���rj��'D�|k����˫RsZ|�`5Z��ocP���Jb��e���2��dޜN�����`@�H�f���l��t�}��҈�C�kES��Ԣ�ܴ�o�������[�M�|2�*��F�r�{��Ƅ
������b���:�� _�/���me<�x�v> ���_(!�v��=��} K8U�Oc�g<�\�����p%�o]��%���P��)A|i@���01����܎�?�����?[����:��!!���,:|��K vݼ��o<��$�5Q3�5�`��23j�}���,u�S��0��,�[�i5��xeߓ�c�i` ��z�����.T�sA�a���Kκ�ϳ.��k ��7�C`"q/�=�Q���|�	L��T��\� �]���D�Y4R[_h֚w������Ê|G���w��~1Cٯ��!������I�5�PV�䣚Oȶ� ��'dW����H�T?��o��"C$��A�Ŏr�;��y�՚ݺ(��)L�sJy��~�N xԡ%ni�'A(���\[�[_��9��`�#��������b��pF<���0i[;h%c33�|.�������C\m�A9��]Z�V��k�U�%��^Bl�$���ά0'�(ڃ��Ր�&���G�j�j�iq�l��#%<��TE��Q�k�$�6�P��ރ��S���.;�7�j��s0�޽��#�p�2.J�
��Y�p�\9圶:��m�D)�(A	�)��������iU�C�������qcՌ��~��#_k�)�!��U���J������|�-Z��/MC��1���$��.��c�����U{�j���T{kV�L�l啲�����_���^���Dzqױ����M��U�� �(�T
عm	��Lq��5��ĵ�V��x��[!�>�FJ��l
6�ww�9������rH����4�:&=�{[@��?�͚��g��#���ȋs^u�F�}�络ʾԙ��H�/s�*�ĭ�?Uڻ��\z^D+|Kmt-�/ҏ��,�|���M��!HD\�Kzs:M�"��{��?'O��6x��)�<�J���_�����B���+�����;&7��r��z���J���P�m3�&���-o� RQ�+���}l ^����8H� ��3f�۟v���m�0Ф�ت�s�[����8�b��+A��q���kGH�?��'�;Q�d]���3Diۋ5b�$wmE��p�	Ţ�C�d������J@T���g��)nRS5�%�H�ca�j>�<�kڬ`ʼ -
�����R�ih�r:#�X|z�s�Eϯ�ks�T�� �L~M�?!��V�z3�b����A��s��1���*��.����QRF�>p,5�]���4B��C�e����L��%=���SX~�`￮p�q��#��B�p�X�p���e���v��X���H4���]��UX��NWII3�,����a�(�w�?)�|��W���]�fR|�`8� #���w����@���%=�O|�'���IXa����_��k�퉀 >�f`��}z��`j�5ت{��:$<b�gmM)x~������շʣ����Ҧ�� �>(m6��R0����2gF3��rT�`�ބ]���yO�o4�o�`�K"#+Y�� E|p�;L��C�ԋ9�/5 �r/���,�P?Y?�����3mv���i3a�O;&7��5����� �><]ѯ��3��{g�?ڂ�rY�|e<�"�s�Sk���c�$5��Px�Qx-r�s���,��[����-:�z���ܷ�M�P�\W����aF��t�-Y�z�t|��_8<KuS��ި@�?|�N�2�����G%��M�'�@�keڛ�0���k �`��+l�P6n�^ml��ޑ=�%n?Y���ث��a�IJ���Q��pinUK�Z�qG�p�Y�~@�|���Fƥ��p�?[��}��n:ѵ����~�����75���<��Uh����<�����;^y��?�C����.N���t��� ި�LI �������_��:΍��|�S0�s��	3�C�+��W�?$���}��k�����gO����9Ɖ0�+���W���頿s�l_,����`Ԡ�xr��Y�C+���_��]�R36 s���PnY��(K�%۵�EeD>��!��Z�N|k'��D��܎�����~�X�%�ih��\������������	}�Q ���߮(�nb�wX	o�R�g;�i���- �`�d� ���<7��(d+"OD	���=����>�Tj �#�!��ҭFf���!W@���'~�_&�w_ؓ���ьp߈7JlC��G O��jb����À`���kc�bp���rԍ��������@� �~e���݂#g|5����w���|���L������R�썃�ġ���j��w���a;��TO��x�]�S���|����%}Zf��T@{Ǐ��f��vۘu��wR����
o]�q9�y:�f(�eb��+J6��N��9��(7M�(4�������?�0�H@j��`��\�~��{K!Z�3�v������a�]�hG�[��ɔW7_�
5�4���"�q�*����p��=���ʝ��ͧ�������w��%ɩ��϶o���ޮ�0Dv�8�����;�~o��_?۵���
�u6���n��<|�K��8���O���~o�E���xq���-�I9��Ϟ>�?&.�&�(����Л_���R���ߖ��?FeĿ_[�j����7W�����n�U�����/���,�?^��{�B�I܏�S�é�7�7�<;@#8��]�mAw����&c��n�.�Υp65���e�j���8(m��Z=��dr��>!Rz��R{;Nz�E�vԳ�ݶl`lu.
#j��b�{pD�l���K$@���/:���@3C%V���,��O�f���hضD��R�u�F���c�~��Rp��[�Z�~�� �{�2G3�W�����?Wa8N�V����y��X�B@@�����m��=[O;SFbT�u��lI �4f�Y�Mp����N:�,��赖.��� *'��2\7��l�m�1	��UK���tb�"�Fˡ��BB8�|�\.+��i���Z�K�w>u(M+8g H����'�7�X[�4���'O���	���E@xk��&�����3[g��3Ϩ��N����
�WLMM)�Q(�p+"g����;j�?ῼ���"��ө�ۧzk�~jw�P�3��E���&�뤥o����^��o��U����3xAA��;�;�o�V>K��|k0pӀ�"<����z١��e݌�'.BZ��n��0)�(VE�tq�˔_�?�p� �Lm��> ;?#ݐc�G9�B�]����xu��G��rM�����|o����˓+N/ޒ%��YgYK~�B��rm�����#o�p|��H�0��I_/�r�|�[������/�)g�v�ʫ,_���&J��܈Z�ﵑ>g�����aP%X�\���g\#��ǈoE���f5|�G�|t�kß��������ԕ�?��+�����eV-^C�V��5�^��s�
�'4S�mG�����^����j�k�k��3tf�
�в�+��meQl��`��IPmZ򬘈���^Y<�\Q�Cm��m��i���"��=�աD�$'�JY/ᩉ+�"���2�3g�U(n�0Rn���d�Ę!al���G��%���e�lr��q�{q�[kSk�`K˦�q�%'+v�Yӎ��T��eտ�k���uo�y�1�E�	��`V<q+*��LY�W�U�-�w0+ˢ׻�_��i�r��=	��堪��v���IgN3�L�����u�6'���=X};�k,�6[�{�ᔊo�r��(Kc�<�a5�Jl�B]ɐP��L46t�VN,P����7ntE+�/���X�\��KL�Y�-lO�lo!(G剪�щ{Fzz�����W����bt秕��q3��
ǰ��#z�����.��9���s���k���(M���޾)�Y�GV�Yֽ:��:��`�m}�\��_�/��X��	�[�����\��	sE"�[�"v4D�ؤ[�:����i����}�]MX�3��Pu\����{Z��:P��ԫ��qy�jtU&�';JZ�se��!������P�`U��wY.���c�
n;�,Ώ{t�	���F��~��`����#)Ïݵ_�f]�L^@�`�l�)�C�u��}"��u`ս}'}_(����sjK���8mI�ଷ0bיhs�v�Ѩ�ĉ��
i=���a�)�.��Q��M�Q��?���.lS�C���`���}�	�Q�y��?�՜YiĀzE�W��뿔�I��L�����jR��}#	�-Js:I��"��Mx��t;h㶡\(x�5Y���jz�=�3E+M�uE��'x������w�E���R���8�/�i�Q.�ϭ:�S=#\�P�������?Ҿ�(c#�L(���@[�^	a�S�Zj�#��;���+>���ڽ��:K�9�}w���a`��	�T�%iz��[@�*�7rC����dʩ��8�x	��@�-�0�9���y�������-��q��QOԖ��d�25�a�k�2���k[��3�u��߯ R��$��7N���r����:�d����g�9���
��B�P�|����f���Z&p[��G�X����z��Њ���������.j��c�\�"�i�!M͇���e�u����0�;��S��ZG�,�-a��2�'����Y�B��Aja�.����Jd��cF,����� �`����[x�ģ/��%�iHD��I���f�nr�(~�&G7�f��̏8�a��&�{?b�Nc����l��F�\�NA^O$����ܠUCj�p�s��l+r�CR=�>���;@����ʆR�� Y{e�
p+���é�g��5i���O�k�j<�@*wZ�_�_؁�R'Z
$!�3��a^a�����<�����f��EC�I��ı��$��FJw[$���sv$�:����'��-ֆ�}�h���ۅށZx���&p��n^��^^HS穿P�펠�Hj	�����̚�(䠏
<C���鍛�Ɗ��o"ѿ�gEE�u�E?g����)������В�ˀ2����1�"�����M)| i�Nuu;I��^@Ԣ�%��g#yS��� ��W1����c��@���B3CJ����">l���b�܎�	�N3I��G*8�鹮"G���(���%�L�f9����&�����ږ�8-SO��\β�vz��dQ��n����'^E�����qG6?p�Q��7&��K����*~�8#3CL:����B[��H�� �&���B�DW�醧��R��NͼK�	�݊ꑣ�����U�?2!��-�
ؼ5��13��Ē�Y�h��׹ˆ�R�]�0zy>QZf������n�&9���ϋ���s�W�{�+���/�L�����
�@�?���K���.�����T�9�8[ee��L�c꿓44*���s���(��W��q�~h�������V(zn�����K(z��Ϸ��n���1���6�oZTN7ko�Ũ���x���^V��^$���\ er�LLV��-M���؂��)����N��ˣEݰ�}�X^K��S����>�]lkכQ%/�>P�R��y���#X�
Q��!¥����a^��L�O�]�R����ǉt��Z���{*+��\����I���;���@_��~÷L�sja�����rV���X	q5w�o���=7�G/�:;i�3
��V���bg:��3~``��Xq ��\G�ݣ�wi6o�~~�}W�<ol��/\�]���=�E�0A�8��+�vs�b6�+ �6�V�uD�F4=��`�!�O���� ��z���}�;����PlA�m����]J��u2��~m-pVx�?b7D�֓��i�K�0i����XU]4��9�l6f�Vx�F��+o��C��/����eϽ(�E`ã�(Pl��mG?��q��x5�����iN�K�Tta�m ��Dk�O�܏V+~�3b]��|pxGH��s���--|�X��#�l��z��$��?��^��������3�UA��^�6ˑP�fO�ʹi�����TS���K�p���։Ȼ,���ϖBɢߥo����{�Ѥ�:O�i$��
u.e�Yc�� ��9�,'�8�oE��N�X̌�r�����J#M�B�qo�Q�5����^�뢑�#9� �J163S�۴�V��|��h�r�^:�3�����o�(�)�-ݔ۳����"��醠��B�L���k�3E�\B:�٥`�ag.����у�
�"a-���8ɟސ?i�*xhs�.�9�o��m�_�1��p�����qaC�{�>��3�z���m�6�t�S���1(��P�=M�2�zrb�g����pV����_��>��ͯ;���:���VvK	���L͗Ⱥ
i�Xز$Ix�vFrb5�@V���W�{}-��x*qJ��9�w[�lϱDFc�4Y3sv�ǖ�c�>�|����CRNb�{,�t.�#wO���)O"�z���e���3��Ux�no�ɟE�,���|�bA,�ه���2�< (/W�F��ɥQ^H��WH�.mA����,,����cuptMe�?�b:ޗ�STj6NzBj0�p[6��9J�us�-L3�`�=��8�q���q�P���g��+��{Fu ?l��ʜ���ǳeı[�>d%	�8�ܞ(|/�� ����T��c?������p�/�4�d��D���5�[��K�d9�`_�q�"p����N��)����]�1��Ϭ��~���C]'zC��c����
�E��`# �01���� ko����e�튁1��������!���;�G����}�(��d���r��*Ū�'�FEz����6�����m3������Yc���:����x�V��t����.��nd֙{�_���I�b�]��8*��0���0�bK0r�C��78�5o��O�0�`�)�Du!�Im)����&�W�1?�A�$�d6��x61q�ms��2�觢��ۧ��E&
3T�V��k=O͔���:K&z�W�(��Ӌ�Hg~(���$�� 8&�pc�����Ii<��o�%[�=�{���U�X>u��Pq�����d�#&�R�O�AN��_ ��!`��I��7^��o�TT��SPR��c1q��q�9M9Y�-ͪ7�U9Q�5�n�Ҩ��
��[�H5ɀ�u~�/�4�b:Τl��C37���< ��@���[d��Y�,s�j٩8�G <��$Uͷs�,O���<4�8�RT口'�:~ѷ�t�"J*���5�2Xlb�?777�M���,8���07l�z���l$��S�������Z�F�D׍�����'D��]��R�ȩ��U���x���%ĵR1?ZS׬&��8�M^U3�����k����f?YG�+��cOj��c�-�\T(�|�l�4���wA��JP~/-1��a8ޘ_�ѵ?��A콊�S�(��P4f�H �'��&W]?�D� �X�'�5
�D�*!:����]E��.�#Р��*���� �,�'��|^]n��噓
C�*.�p�u��x�V�?����hj=*l�Դ�G��ѵ��COz����?]�_�oV��%�g���i�n@m�Ԟ;G͌Z��V��εkJ��M8v Z�ɟܣT컧��c��_��Q0<mB��_�ZSQ֘�?���N
B����M H�7�` �C���wW_���R��	O�nK"R�;vp:
Ѩ�m����Y�<g�Fb��-���4����{D4�f�[>G�gRT�������v���uf(�Pi�ųc��6�[nT5W���J���}ц\��86�vīKD�O�7��QǣcD�E��ˈx{���3؊���4�sqHt|�36��B��Y8 9?�f��?m���:]�m�D�Q� i'�S\��]�?�~�hc墵L G��5��X�v�8۲>JCZ���d��~Yׯ��6�n&�,��qMG���1����2�RX��׎\J`y_t �� �p|�i�#`̲��8!p��*���Z��;�ʺ�c��\�_��1$�V��B�iV�����?�9�f���\0���ɜ'�,}ɲE"���_���L��D�ّ���K3S�DfH�⏊b�+����鐌U ���f��L�����N��N����u�O~x��ߣ��e0, ��y��[����v-		*��!�Jq57�e���B�o������6������n+�y��VItf��$��g����Oq��!�z�����{ͯ���@��*�6(�~�n�D�~r�����*�I�?�X�6�6�J$ �y\o�z.5SV��	=�f)ݦg�
���)����"�yIU9���A� V�cQ��UM�>�eI�NC>a��
����F!Ȟ��F�g��]m`S
=C��*���eQdZ�h���_�l�(<�7wΙ��Ű���P���1��C��\�}�m�:�u&2�+YȎ��VL	��Tw�����i݇�̻^-X=߁�;��7с����A=�#P#e�]��ȏ3dD�;#�ϙ��88'�|��?ϧ�:������Q���Bk{m�����D��y=Y���~��'2β�����Tcu��O�a��u�F�֡��mQ1f�(3�S���{G8T&μXx�!�H��si�X;r�q�d��S�w��>�z
��Q�Ԧ���85�Q�qj_Y��2����1�p�����w"�WȗˮOK=�'�w�+�Z�YN��rHݬ:���~���M&r�7�؍�?qP}�� �Y����J�y�Vf��fs��E��ݍ�%Y����T�?�����4����T�mUj$�ۗͮ�O'%ze�4d���v�ɞ�~^9+��ji�)He��>n��Y��u�xz�~���{�{�`�+%��m�7��?S�ô�I���tY9Q�_u�#�}�K���CZƟS����W�&���^X�,�����1e�-� }L�!�qt.�Ҟ�; ��/k��{oU�Ǎ)%T*��T�I{�$#�!ٲ�;Q��d)�}gȾ3e+�:��0���/�}F�������s�uuՙ9s�����|�s�}f_�q׼�S�^{u=�idL��Z�V^nn���Q�ִ⛯p34L+�?�k0�e�o3��THm���hgX96� g�w"���ﱱSkN�<��#�[�̡�{@ �q��?S�j��ƞ� � ]���7�N���eXJK#�gT���hJ}A��X���}?j �����2��{���l�Ŧ��-u\Y��b���Wʋ}�6;H$2˼6�{����N�Ujf��<�zU���N�'�\�ۑ� �	;���N��ϥ��|���\o4^Ƅf瘛^S�IW�ة��yIݙtޟ��F"��C8\��p(��/��B���>��L��y���;��n+�� �^C���F��j�����	���6+z�t�O�(cP)7��[����I5'0H��Cw��t�FGj�J��|�Q_@���.�{��q�R�� -�bg�WNJזI#߈�u�$>'K[��U��]��W>wJ���S�v���\�kǄ=�⥟�)@�C��[Sr�;w<G��j�*��I��z�D��L[��#�c�|�"������N��u\.�6�hc����:����kB�����9MT����1Y�iת�[+���v�����;�T#2}5����(f�����_����4�9��Y�]�����y%nߪkK�X�vpE���cH��hNi�Xe���s�d��`���a�z k5���� ���
�e�ǳ;;\���%��S��(�_�H|���	���Sͭ��:"�$�x�=�������E�;w�3��\*��]f\�����ajs������9��zck�l;�v�44�Ez+��<�4��f�:ڦ��t�ѳB??��i5�x��h`�*�V5�@t��������\a9Y|
����a�kDռ7�i�h�3ȖQ�L�"��p]���f���i
�z�C�e�ӫX164no7e��$|���[�9U �uv�C���U�O�.!�(���IK<��x۫��9X�#��`�w��J��cr@<�ӐXwK��K���z �Ռ'-����\Ҟ!Sϗ-X��UZ��g���Z�t.�]��$���'�e��rLI�9����Lj9�zy�E�c䴅I9b`d��d}��R�m����{�M:���v�-��/�h2F���F[x]^��N7"nv o���'��^��|�ҕ�#�4��o<�)�O��'nO�����M���q��ݽ��/�Z���^��{����s,�������R�Ʋ�� �k�����e�-��ˍ�j4'+�]O-,�;\����c�֎_��>�"p�;_���Z�u�g��N-.��7�����8+�
Y,�k���s�<8�yN.1�5�&8�j��ƀ��oY�62:�<I\,G����i�E5�
c^�����I��&�T�%L�Y��G�W��N��
�	�Vrh�<����z�J��.磔�0tK%���\�lE�0�K\7��'Z�]�ix'�mz��d
]h��!�N�%�PMC�9\��:��@qJF�׾�K�p���b�%Y�<�A1�}t����;��ҝ�����D�q�5i�մ�;�3zH���"�
�R�Y�iv��&�c/C�٣����-܄�Np�P�y�Y��B�L=$�!_L�T�v���Q1��\T4��G��sY�W["�,��Y��W=�� no����70�m��GO��k�2��3�^ǽU-�-�1~� �3��*�!;u�d�RG�)��FM��������6���Z����}����a�GB�&�,>��ӓxk׎�l���hY8q����(P�̼ ��Bی�egR093~�(&[��ekrZ7��}��d?�]�ه]/�g�9�Z�,Ʊs������i�
���A5�6���45#n���H������p�@��44��Q���'���L%=��˟��Ar�E���Ф��T���u��Єڢ�7J���[~P`R�X�ʺN��I�������?W`0�ſ}��}�a $�o�ԛ�����Q�豫������P_᫇��-��e�4�$U�n�Ӫ��pn�.�����h��9��6�0��JCv)m�?�@���;�	��o��%d���kwk.���̨Fg%�����qh���yR���1.%s�k||HK0�������Q�u�j14��YfoWz�r�f�����ۋՎehh��0�#A���y���\�R�ݣ�f�8��˷4w����C�'#�?�C��黌�c��O���֋���솵�<�����ku��-�F���z�0��_M�-6�&a��!�ͬՁ�&�Q�@6x�͙~�͛*h��$��u&����|������g�����g�CO	$���2�h�]2�<�t�qLA�!z�#}] L���O��tN큪"�w4��Rx׸*�Ё<���+<7�K�n��(:a堧	 \�מ9�i�lee�JM�:~��z#�Y���y��wOڛ�J{q���q���N�+��*�#A��^>���<�y�їkh���~m�~mx�-VMS(LGNS��gRTX�cLE�e$[60(���ݠWh�Q^Ն�-�ǃɦ����tM�����OAQ�2�v\8CZj��A�"=v�Y�u�����˜���~Sj�F�~� �գC�m�d����$3m��P#�M_ZB�2�>p�lW_�"�.�Q��7�0��wĄ<aON:����z[9�*�<F����m�ھ�$3L�*�U�B.i#���$~�h���6QͰę^�`(�[?�����A?��׸����-Il�]J�[�\�iXS-���}�JT�ڱ�FF`�R�$�\eѧ�欉dj����y�G�r��j�ߴ/��Ὦ\ ��B��$Djq��R@!��2+))9�r\[8̮�3�����(Cd��4�O�oB�9�`}�ϖ�t���JP��k�TO���_�l����������0����B��6���:7�׋v�'�sk[�������PߤZ�jp��]�3,��[E��Ї�Gg����x��&�j6k&T�QM�l�$U�V���Un�N�ΙE���o��=����"�������VX
��m��"w�th����۱0��Kw>`�0���GU��k�Q7c���4t�I�<�w0�԰�1��[E��W�h��F�����i�A���'��Lj����͡�s��Ù��Q���]e��[\����=�,o��-��IPb7�.�c9Uh}�)6�2��Y���sܮ�#�u�5*� �-�L�`ee�^P��m����}��V߆�8?�#��Z.�9L� 9)���R��JAc2^��
a-��"�`75RA#�ZCN�4���:� �=OS�"�F���Xښd�͍��`��g� �7J����r�:��OK�o�*I�Κ�y� �c<y���^ͦ�,Z<���*3�?n��/L��ɻ���e��:�`"�����V
�rˑ����*L��5Y�y$�ء�g�y>l^�4|w^���[�a�/��SM8��pV�ϻ`���4�B�8��t<x��j���0ZYhƿP�!�K��b�������(�;MZ�����)���w��2�w���4���]�r�}�I�\�톉���i~�	r)cyqڰ��g#r�|��(�������G���s�L�u*�� ��tFJ��b����J��}?4��^����#�Y}��Ι"��dW
'I�+.R~��"��̿ǜO���%sRwę�ǁڏ�RwyR;� �%u����W_�`�,�
PaZ�\���.�饢�� �LT�E����I���fJ���j��q���E�4[�_���U<�G8�A܊ۛW�@��I��<[�8���M�����|�~�K����Ly& �0-���-?�f�+�Y����9�Ff�[s���Ee=�o햧��:aD��,��B"�"�K,�F
�;<��xX��Dp��&�^�MS�;e���'��y�����A�8<]ֶ6��Cq�S4k�~�b{[85��U4�|��7�r<8t"5�	�Y\5N���l�n���@�]�o��!|L�#����z;D�-į h��Y�!���,�����n�٬�YH/Ú�F<@�)-0Hs"/eY�c���q.�����;�����H�Ռ�sc5�Ɍ�����c����<������|s�7�}�q#�'N�n�*���!�[�l�:&��ς�D����ܪ��j�Cgt�ڂ&&VZ���? c2�^��ոWl}/��Cdk��#�s�@�L�[��쾇Xb�q�.L�
���C��fʖ���Ѭ�"��|s͞V��peW�BwW�k�3U
�������[w�zO�N��_Vӳ�gEVf�A��>oٝ�K3X������g��D���:����� �7��}uw�,�ҧ<Ǵ<�qA|_Cڌ��N�������)L��Z��������C����4z�?ݓ;O.�0���lL�@���ή�ܨˇ5b�_쾶�-b�g3�?l��?0�&:������o�=��l�T�Ev:��;��;�	��*IV��TK?��֧z�7�*Y��B�ᦇ�AS*��0#�ZZ﹞�H4޲5T�d�� �ދ����O��<��,x]��6���~	3>���}?`���+?6Rua�K��)�?��?7�ߎs��"y���h�T>\=߁���8�i7i<��|�"��� �B����������~����V4�����s^&�AnX�Ț��R�0>�o�	�nV�%��P�Ȓ�,Ȧ�����$��8�c�g��d���J�+��z��W볚���,�GU�4-���,��z��I�����WK���6dO�^4�[J�l�{1	������W�$��o�e��[��n�.�z�ٙ��h�f��F|-8ۖڈ4J���������M���KP�=3�4~���N?f^���8�0I�wvψ�QY�$O.S�M��q��Z�K�K[w�K91ocM�����4���Tv�X�Z��;B����XA���3[ ���^�q{V/r|i����Y�\# 4-{V�bnU�a�O..��UԚ�t���:hVL"���i��!�P��Xǀ���1�SV�_W#Մ�K2���*�O�X���loY����eY��� +-���*؏���#�*�nϖT���g$�>��<h��C�/�\��YGg�P�-+��YY�s ���m�ӷ;� ~\?��~�	^ �7ESLa	[�s�~���/ڡh�ۮ9�Y�]��$ �Ύŧ��A�+���5�G]�P���"�qr��W\����>w]��Ȅ��#�*����/Pkv�/^��2v$�歝Z
��O"h�q�o5��J�$_��{�̈�s'���@v�����y1h�iɭ`~� ��t=���|hU=����<�[ֻD�K�'� W^>PS��+��l�xh�9C�vb)����T	mE Pscy6*.L}l���=���oq�ߝO;$�����P�c�������Hv+
OM?9�nj�c!�u�4U���Iʾ?�5�cêk�͢�m�dv}c�B^F�)�b�YE�=��&Y Ǫ�h;J��F<���� P���)e)�x4�4�e�Y����<��=9ʍ����U/)�y�1��K�P7���9��G������2��q\���<[h=,�־�D��kr�կu��xM]�5]��Ź'�Q��@�ڹ�[ ��o�㚛����P�Rz���/$��;4�p���2W�]Ci����@o�k�X��5�Pɝ��j�/[�2��o��,_�Z"�f�=l�����J��_�*h��è=v�+O,0���Q��c� 1/��:0X�eˣ��2�6�6�j7�s��^v�a tE����+��Ӥd+�4�i}�x���r~Ԧ2�\��-`l�Q��ve���@���[|G�/�K��� ww��u��
D|n�v�'�|t������ �Tx������p��i6�� }��k�ʢ�y���y�]����7ې�w����3G� �8̙�rR���BUE���Q `'�M����%j���W�Y���ym�����%��h�)u�L��ے�谝)TI�x��� ս���Di;3�`�O���f���� ���#��&������rZ�� Xj�<Фf�����
��Z�Xy��0�痓����Y����I	���1���r�^܃�pk@/R�_Wl�v������M�К��W���I���_i��yc�X�_�x�k7�Z����(h��&2@�-��.b�f��1n���:Q��@�����Ԩ��b뚃�����mC�wԶ�Y�:�b����s��a<V�.f+t��#:��3'�x s�,C1�RjH�'C��O@K1~.�*-��@����o}��v�;�ԛ ��ښ)bQ=��:� �r��*�y�䷛���J��l7vL�![��%��EO ��Oyet�	Y%�Og�5�\k-�<��2=9�Q��Q|�$I��)����^�&��qN��Y4���!�M�y����� �T�(�	���`'�l�邆�;\QZ��
z��a^عC����$Tc�ŕ�]�T�RB��ؠ���d�CzL1`_��Ӌ��A���GO}G��0�a��%G�gz�J��S��1@�Y�����oy,�⊢�R&UM:��gM�mQ�'n<�`�5F|��Ō�Yn�
hxꤤ��-���tl�մ <�=?���7!��1�ֺ6p���H{��R|�˕1�L�0wk�|'w�N�G�����5��沽 }�%f����'���?D�zxj�Y�|@�#�4�Tpz"�6DM��5�Z辅���B��j�3^.�~���G��5�h�
��w;Ў&.��i�eo�9P<�a��ſػF�^�K����r}ĉ���>G:
�Q�K��B5�i �Y���MÜ�W2�k�*c:FX���:��#��3a�yv{��H��_��5#��7e��$De���M�O��.v_�=��a-x2,)�D��M�4D5�������z���,��:
DWC��GRr�-�P�>rl��f�9xX��P����r��]�ـ�z ��VֈzT�����C��<���[�? #<�T�����VK����QX
E�@�]0�(�Z��'[MC7@)&d�Nww�t7\�$�wdK��j�d�~�g}���w5�"�cx���3�[�Ά�T��q<oÁ%�Q~,�c�1#-*%��3#���	�z��,�.|3B/�W~ѕ�6E�%C�Z�{	E�)�v��f��n{Aap8�&D��G�  -1�u\_�`��b�xP�^�6	�e|��0,�O�y
��_|�����x��0��<�b�.0�4�ZBҀ]/���j�ݵsj����l��T�T�_9�@ᓭE���4�pq�I�eXȂ'2�3�&0t�6>�:�\��5��B��$瞮8���'� ?z;��F��ڂ6A���
�S�DK|��+�fB�f}C�v��AW� �'�q��-��#$h3"Z�z��E@�W���O����x��6͸�Y����m������z���f�pec��&��Ł�f���9���V@�1 :��F{�[E|*>	�eh�8w9�	��X1t�' �N���TYoW�I�|�W&�-8�4�.�q�룠�����A]|�H_��C�y�5�^A�Aey������	rץ�~PV����ŀ-�Y������p�����('����B3��:`#T���c :A�ud�i����Aj�k���Z�dO|�}/@wJ�5�rHp�sa�=�#DBm��$X*O	v��ͥ��ޒY�$�{������@����֐�⏑*��1���^�1��	��CE���F m�\K����K�K^�G��)��i!̎ ��T��wX-���2n�~��H�y����\�����ez�S?��͎�V���;"1�
����D�p�H�d�nu���k�;r�	
���X%��4�J7ᢊ��R�m. �x�2b���x�^��H����ji�]���M�!�����t��QN ���a�O݀BU�1Y)�����!������:�����w��P�Y�'?�*-�pY����x(�v��DAf�.������nx����ݵB��q�]���4�&�~�/��߰�������<��1�#-A:�0t�@%i�  ,��� lњd�%�I�U��<Cy����)������S5;kc�z�����?QrsCϿ͗B{�#�Ɩ�J*���:i��#c^.�t���K��V��4I�-W�m@I��f2D>Tj'`�����a¥����	x@"`dxR�"dԓ�wg�a��F��15}ֱ[�;�e���7ӫ+�L� ��k�P Ym��>��:P���xoM�<�%U��zf�Z�>�9�+��]q��'��>R�ٺ�k=�ꬖ�f����j���Va�k�^,�L�@�=42�
���+_���hvoe>�Z��M[���:UD���1�
�����oЌJ�j<G����7� 2 �3��7Кɼ�&[\�6�_�SXC�($�$D���J �,�f͟��l�8�?�杨����z!-)�j�4�AB�	�=0|��$�F��V�����/i@=f�U�Ý���Co��*�2:QQ�|9�e�GK儊Ņs-X�L��UMb�����>�@�-}4m�I���JiA� ��b�cۉ�A�������5�Į����x�e�aa�����cN�˷�0蠟h�0L�:u����o(����N�n�uw���� D�D��;���<���R%��J4�!G�o~�}e��$ؠ�Lq$~�S]8�df
'un��Yy���e>�+�"*�m��wS��k1��Y ��^�����>�x�}���vj|^Y��N��*Vn�n�>�/ӧ�.�ngno%U���-)|���q_3om��/{x�[R�	s��U�6Z��J�a��.6~$���:[�\����"%z�`�������P鋖�����_9��9@k7ɝ=1�B+�$N��닥�h^���E�[`}�����ל�4�>cu[�:	�<;1R���$�^�M�D)mG�\ �yA��!�PeP��Б��@��T�S`VrƍZ�5[�\�4���h	��B�ĺ�J���:�YѪ��m���B޼8g/��!��6m��D;�WJ_p����:�W�@|�<G���g�Zϟ)GJ﬒��ά0I`k���������{����lm�D���b�v���p��.�Y�g1��O;oq�0��?QZ���9�3�{���L&�^�=����t:/���7՚��Κǖ�I��绬����ŉ�������E�}��@��F��HP��}���}a%�{�Fs�u7��1$���V��LL�r�z5>4^X�nAWà����F�3ۡ�%�\�f^��mv=w�KJ"Ag��B!b��
S-7V���v�N8�H���ף��3�@�Y#B ��x����j�-����۹]Z��U㝶�"],ݡ���Ա;��� �@o��%�w���B W��`ڮ�=WEYP�P���a����(q'��@��Ύ�ó��{���K���O�G��am��J���:{�VM�E�g-u�n�9�[Ϯ�V��N[/��s9�a����X��V�P��Z�0�M%#��U�:�ɥ����G -�P�	�lg�&�Q4~�o<��U������P�����6���d�WY<l��*��EFpIK7�%�$T�"-�̢����Z�q����bF{D06W��Y^n���_�� ��B�"�j��SV%�d����ę;?X��U�V���\��T����T@çӐpw�c������B�V�ft^�u^�UxcT�V8���S�C>0T�u�O��tk���o5�U��}R���9n'�,X�'��*���l��t���ם��.�G�f�l��'׃��G`�I���:v�Mc-qj7�ɻ:���BXo��'6������J�Mu��ۮ,���5�Q����1j\~�Sh�t���-�k�Zp���G])s�L��E!�����{!Y\�[;�����%�_=�M�p�������[xwj`�Z����0�������}�:�K���xj:�tuQw\Ra������w#�z\�>����rS��H��&o��@akGG�M�+?c:ta�Q�*�VS��4��}���=7=�d�@@B�����9}���K(���7���B_�b�GxGn�BՉ�\W^ |�N��+mjI��
h��"/�:wupݖ�{
3%o�sr�[sU3/D��G��f�C/~�=΂[�`���/�4�_Pt<� h�]khG��#�(5
�B�]�u��0�\�f��^���u���5���`�h^�ur���%��mR]�/D3�]���	Ny��WALS*������_=�˂���;	(�&�H�	 �M��z�3���_'k^�td�.�-���I<D �a9�a�ζtN7ov{���C�J�F_�O{�>�C4閣��P�p*�>����z���J�^o��5"���T;1-�u���z��vXQ~�`̓웷�m������W�R�P`����D��n�g!���2���m����!�ͭ�����"�j8Dom)��)��%:�폷�əQ�G2���yp����������f|����`���d(�-��6Zm�]�V�f�5	��ef�:��K-Rq^�̨�:v��̃?�g�$z��A���q�OФP��i�_�;�&�.���%���
��*�qѪ�>��d���&Ce��L�����ǨV����)���U2�)z����oM��(���1������,�8v$��D�WUd���̮_���$
�@� b�ʡ�?�B@ m|����~m�>%Et]E��Pk(��r�i�b��uh���
���;�8D�}&(� ��J?�)~���~_��Pڥ���_�\,0?��7�:�x��o��E`���A���MT�YĚ���&���N"����D�\�`/��yvz���9���o+򸛊D����3^����ƞ���bq�z��5<fz�L�Y��*�7-�2;υv9�����A~�:{��Q`=��݅;T%ӱZW;�ᥠ�VЛ� 9ZD�,s��?Ġi~��sC�B����\*�d�l-��W��Dorڬ7
�+��+��7��֯�&���x�UY��{'ʨ"仄�r��˚�'����"3�⡠��[�ꬆl��t�O?�;�S�*z�G⁼��> ��Xc��]���F����'�_B����߶;�DTT����d��Ddv��q��co������a�<Q���۴��	ǅl����T
�o�^�k�;N?��w��5jb��&4��*'o+��[u�K|M��Ё���'�]CzG��K����c����%�&g������&��;�� �n�����hRayK�������=C�X����W�a���KV��gF4>�����۰'���bz J����"��&oN�j`���!�kU����wWA�#�H�)&I��o���mmٺjĆ���K��K�L�M6�=@�J��z
:�0�]q;�s��:QR������^���?���A�Cf��yHx��]�Z����Am�pg��J�U4ua��o/���|6�%�����K���}���\ A��X�F���E��[{��	�&wf�o�2�S=0�yE_h�oXx<�<��Fn�Z���1��#qo�-N�����8v�C�iF뼘m����E�g��6�4�AIBN/A�Bw�g*�l�`�����ݶ�k�@ID��&M��5h�Nb�k�'�!WQ�p�c:���S�w���T���E|b�J}<
�>G��~��t���G&� ܼU Li~pxmrN�;�`���8���cFn��m_<I�k�k��mOJU	7����`��1/� ���ˆ�ET��w�x!xӤ���ó2��6\#�}X���5��/6�ʤ�������N����,��T�bn"[�L��f��~�m:��W�p�I�PT{?:-������ ��]"C�H���[*�V�F·����U3�+C�q?�Y�^����y���j�{:ʞ��[G��>��%#��`�X�����|m��&H�HL�/ߢ=�,^%�np�f�C�NOQ�t:#1@y\eo:��6(����H%V辖?~MH�v��
Q�fnɊ���xPL�_����P�J1i����'a�rW)���<��",����/H�������Dn ����|j"0;J�zN	��%�@k���)R��y�&���CGni%�l�����&�蹾��۫�:�]F¡sꁐ�]�6��5����`�/�K�\:?���p�> }[�'��R)?�
�\泰
2ou�����B�l�W:��b�U�c3���h���1\\S�N��1�^a���~؎��ؽ}�Rq^#���,R�A�Ӝwϖ6�;��!�Rp�����H/�\�f��,P�<�4n5��� ?�7�ǮtAw]����1�j�)��tzh�4t��F��`rfM�)����������[Y���<����췕؇�mkF0�O�s._�7Q}�A���c����\�f-3�
m[�nn�_U|D9�	�(Wz�0_ z�N2�:��ؕ�΂��X�=2y� 1~1��Tj�3U�>u>4��7am ��6(�B��>��O�&N-������>t�P��QM�a(Ѱ��8qC�+�<8���h�eli@S��O4A+&����|໠����f�*>o��S�$#A�<$���)~��s3I�f�ږS�H�^���c�#��Lh9�r��6����0�P�]�8Ӄ#�ax*���)gǝ�g7���R$�?(tn� �P�!�w�T�PJ��]���6i����.���������τLM��U�ܑKvk����K���s��#�:�>8�j�v/}�S,�ϗ�H�B�Ø��@�^K���y���7�v�zO�$��):#�����ywV��d�\�9���y�/ӵ!�sbDU� ����S��A�����ӗ+�{������GH�6��ӭ��W$RLg����5'�>�$+��r��r4v+'��٦�U�!lD �Zu���}'��7�7�ٖw�;ee���cF_H� #Y�"�0�\���)=Ⱥɸ�6�RR�m]�A+�#��E�O�0^^jn��I�]���_ĭ��ʄ7�"З@��>m��f!��R{m�t��w��Y�N���'����a��,�(�ǫ��g�4���-�s\p�u�GҲt�i�4ҷ׺}{����U��TsV��[]J(�S�aN�@�q��J�}w����E���U�~�/�(��n��˼�L�a�DRw�p��������C���΂���KMi.k��m��>�
��eOW.o�㾘�E~r#�@{�D�v��=���Q�$L�+��1lS$����83�!�}��6ƌAP�L�B+/�T����3+(�S��:������-?�/�<o{����w�z6	^����DRg��c�s^�D�r�Bn_��c�� =��[4���qN�ob��%��noG�-�/�@�Q�;,�9�
��)�תb6G~�H�D��NH��Ylm|�%#�%�n�o��%�����r:�^�j=pߓ�΂�W�$�BJO�)>!����G��wV�����MЬ%m
h2F��s����=F|�vrw���vݴ�i]2j^��[e��|�k��'j����� �)��2ԝ�M]�)"px$(*D{�Xx3�����|��|@�`�����d�٩z��3�Λ�M�����O����n���׽xIU�?�z�������ȩS�r=�����N&���"�=_=�t����+&�a2����?_��D!����x6w�ծ��0�{���;v�0��'�CY�fϮ���ջ�\�͜��x��<�j��p�L^yf�������i�*>'s���xY��l��%����^q������*(���F���X'zO<�~�r���|�F+�~��.xMg�f�0�0n�iq�?D�����M+ڣ5}#��#꒙�+�R�Ě�}��ϴ�1���'�:��	2�j&�]�;<Qt�S�k79͙H�~�}aey�a�.����ԫ	���D?o�"?��cV��x9nO�����1pn�ؽ�<��*[���������[����n��{Gg�F�*�:!�Gw���C9���s�N�>_���h�K�k����ѓ���&�w��|(y�P�C^A~;d��	@D��搢p�}��Fd4�G��-�����d�+d��[�&��{z8��W�/��gJ̼H06=�v�,{=��}�~G�#��>�X��DƸ}�,>�\�d�>���M.R��'���߈��Q�(E��èoxIݧ�*0L���dҴ�_��It�u|�V�,�g��::���tW>��e�O��^ 3c�Gr��&A���{=���*���g��C .sؕN����kP�K�MK{v�/�*4Iz�a����<He��b����y���l`&}�w�![4<�"^O�ODa`�{�3C���ny�@%��[�>�����C8u�4n�u.�/��p�u�w�1y�݄K:��ܓ��"��C�um�a�b�� �]A��� ���,��D^�3�@u���ޔ=2;��ܟIC�0{�M�Nu���s=��k�g��~t��|��F�^ty�O<��/�ۯ�z�x�Lf^�M���wm��S�E��5po�Ǩ���]̵W쎌��7
Pҳ|`𚂂�^ubN��D(�9���ͼW��ϯ�~|}v���`��܇z���0���dcP١���
�,4�L��>o�u�ac_�sz�_�]^s���:����υ�L�E�#`�'�J�cz{cSԑ�sӟm���0��ד��Y��{��x�r�^�H7�o� �}翗l5����(�����4�*s_d��}{{�d��E��E�N��x�9� ��Px/���A��t�q˲)q*�8�WY��n��q����y��;��̜̾9Ň�E�p?��g��ㅕo���#����{��ͥ��-� �X!��k������i��<?��6��B�ŷ!`���g�r��*'p��a��:@�&�;j���r{�] ���s�=�7�NV��Wp=��
�'��ӊxI���>���,�l���+��u$�p�i���{-c|G�fPPWP�Ox��}Z�P�M5�����Y0�[W��{5��=��Io��	�!�߇�y ���A��N��-=�O\�z�	o����u�o�g�i�x}�Z���+��Y�TO��@��u�6���3fR�|N���w�_�6�y�J�r�S��um��__� ���ٛRy �Xa�����I�l1M���Hj�UW�r��>�>P���PV���;�#iuѧv/�Ds I%}V꛾��H��5+�7���^J���+=�q��~�p�q�MM�W� �8��>�U���-<l�)nP8��}9�!ea��k�e��L@�ۣ�"�%_C@Pa<�#�%)|k���ly�����^��/tN+P�W�@�X��-D�^��S���%���9Z`��t�g~w>��2;���I{��Gb�Ki�E*���|�\5W93��}L���z'<����WZ��V�#����O�+-���oޫ.;��s�.����&{�����K-r��>��8�Ʀ��|jݎ��ϩo��m6�x8�~[��W_j���+"�����������3����(�Q�fN�{S�^��K-V �ޤ���ǔ��0Z�>n�R�3�����A�D���?`{O����A�~o��A!�������)�<w(U+w�?�7QV_��p͚�&���TC�`��2��� �޽p�:^��m�\�3�WXT��>ޭn��i���uh�* pUa��w�@��p�����IY�y�jGg�}��4Ҹl�Ⱦ�r�Z�L��kj
�j���9`�"[#�^�ϑ��5}6|o�}q_ڠ���2HG�|�Qާ'��-U�e�Z�̽}_�_�Tl���g$�/�>�^����%�3��ISضqا`!�;���*�|{�5#����	:�S��#��b���H��/D�_@d�9
�o'���rxϛ������{N��,�3+D[��Q��]	���ꋀ��)�M�o�S��N�����l��dC��nչn������b���[��5¥C�'�ah�nv���	� 7v���,��	�����7���t�����_[ YS��7���q��ޓ��;�w����ѿ�G����;�_>�W�.�}/��Kr�;�w����ѿ�G����>��:d������삥��c��bc�n<���NӐ�&g�pq�KK�Q���K9�<���ڒEG�⶿M�� !�ꧤ�'~r�|a��x����KI��钨ە�ݮt3Gnp�m����^z�7����K���mPT��r�}�d��2t���=v��*{U��Ap�Þ#�����?j�S���ߔ���7�)�M�o�S���ߔ��)_����g�M�G��oj���N��g�t�R�}?阉��;7����uG�׌}���Ds���r^nU�ؖ�`������,�)?��˧��a��|5Q+�ß�{��8�m�����?Du��b8
�c�M
�
j3^��(Upkt�ޞJ�9֋�iz����ogP��ol4��)(�����;�9����:�=��W��g��YyO<ja!6iKi<�e�]V�Ս)i��,sg95�/��������5fސD�ڞY:��(�7���_W_�&�415�k�f[�i��n;�Xx�UG�?M�� 0_ś�fw�7�\57�R�_n���'�%6��E���YOŌ7W��d��3��Db��^ν��j��9>؀�
����f<�X3����%��X��b��g�� "$RL�SH�wTK�Q����?p�|�5����������]M$-t�ǥ�ZHz�_<:����W$����ʝ�%f��ԫ�o�%�jNXwq����k(��qp&j���8{$�a�ps�Th��$Ĺ�H��G��r�Ֆ��iq�{��E[-���'����<Z��f��U�!�a��T?<�8�̜as��)��cǎD�sM%�&���b�����L�V9�;�����$��"�V���>��Q���f��Q��	.($�Oo���͵���؝���,VcM�۸o�o"ی�VX�czg����о7e�ξuُ����f�E�`9���]Gq�>��aN�-FZ��3 ��4��8�Hhc�)['m2:y�%�mT�d��u���q+�	��z�O�S��}qH3r+�ܶ���-�pu}��z�1:�СIm���?��=���j䯙Pg9��^������{�%:�IKTg�e2�F������ԛ�iWu��-a{�m+2-PnWn��	٪X�-ߺ-�S�������1)��n[��[߳�mf���MƎ�>�l۸��r�9W8k�F�?L}�J#i�e�eᰏf�zMb,��P��[�飽�7���둑B&�o^~�L���Z�N��ά��v{��T��k͊�K��&���{i���_N(�����1����z��Kn��1c�y?��\��BYw�%��ޅ`�=���3���*�ө�y��Wfr��g�:T�5�n����fI�|q��r_6�_�ܡu�`�i���Q�[\����/��J�@{�,1�57�Tm���R�w�C�.�
++��<ΰ�\y=��.�Ƙ_��r�ڊE�{7�կ|�����A+��"0���+!�:��Io"���)��h���b�3�	K�(zS>\<��
���ŝ��|�嵡�����3}ȥm�LVRl+8˝�Ě�(g1���Zל�%vC��w��W�;����7j�c����8����k;���>�M	��iV���#Q�St��ҕ�#o����q�q 0S�ɦ�o��A����=c��@��;���ݽb���
���O�=b���+c:��iV'F�(n\ǧ�%�/����q�<o(�C����U'�MƎ��[T&b�EU?�عf3kt�t��d��j���Ғo��ƌ@��H�r���sGc��e̓�+5h%[q�?��i�G�ګ��ҫ��3|UUx�R[^���,ǵ���:̾>#�RWR�f���'CzG6$������l�\ΆN��G�M�úu"�������JW#��5�ւcǅ�'��j����c�6�����7���O��dJ�-�{
yAH���������?ԽwTSi>ꌟ�,���f�(Uz��.���;F$t��"5
қ�;�K���Бމ&t!� !�s�03���u����Z�i�y�w�g?�>���`������Xxt����=�eР�SO�d�'K�"��o��<5kk+�ß��4�`���Մ��	�ZVah������(������a� ��m�tNx�f���+�Y2��Ӕ#,^�������V�j=��-D�$R
��Ï^G'PL��� ��ǵ�Ҵ���(���'L��������ܤL�'ac�u�"{zz����	�Q�Ͱ4���^��, �!�\�8�t�qN��|�XQBG��/���z�������璐r�+{#�Q����F6ܧ�� 6��i_��%�����ĕ���>�f c�O����X�pR;�އ=�
�?��,�h���v����L�,��~d��D�>���"�#�U-���s�[{追�~�\~�U�����y���^2�20/��%cK�Q���m�|����W��_�I��f*�B-%�]�c�~|WVV�K�W.G�R<K/�c8Q
���ܝ2����Q Y�&���-�F��ԏ8oC�
�.��^j��04qWG�7�s~ Lݽ�C[Q|�������xzTw���Ķ_�߶ �!���!�4���A�7�����s�ec�����w��'0=i�t�{��R�|�[�q~k�������+���U����:C�Y��/ɴ��@K=��w�hU��F��BXZ�57�X�aЉ��CIU� T� "<���u���PIz�l��RR"|���P���7��#�N륿 B�]�'M��o�7tg���������Tm xV��v��7�j/&{��'i�I�p7az�(��P��!��E�^e'�N �r0-�X�G1�\j�}�}�d�))2A�V�xq��.�����*�A|9�"�O��&{�W�笝�-ur5۫5��O}��s����B3�P�0T=nڸ���� ˽�jd��b�4���"�@~u1�.����D��UTUz���W���B"ha�U�̦�yu�ӹ�͓c9�2zCd�ԖR�K�ʟ�a����e06�w&�G�(kw���EW�� wb�/k�S7Kqk���������8����,�1�����ϠQ��$��o��4{��o��/�=��=xŔ�sU���r����¼*�6"t-��4��tTo9���!�Q�,B��o�Iڣw���u���N�7<g�g�;� �Y~X�x�H�?��(�/�˸	�4D�'�i���h0#�	��*��<�JQ�zoٵ��Q����;lܮ�RA���g�8ҍ;(rE%e೨�c��}�G����&�(wj#��m���A���w��͒����dUG+�s�8�$Mj����+q��wܧt�	V��M�I��lh��R,��K%�Ļ�ڀ�E��W��{�d�Ǿ�]"J���5����0P�V.n�eal��Q]ߵw�Ta��DǴ���3(�ٰ&�%e��u��^U\8����2��IR���Q<4��X����3O>K���I%Wl�1���[8ք��8�k�w�I���w#o�
�^���9L�<�_��������߾�'���B��C7�E�逥��"���{}���6�K=��kr�)��K�;%�Τ����z�� ז�-��}3&.�~;͏'f ,�C6/"�>x�����:��?zd���e�o3M)]�������ҙ��Qޘjt�Nl��`̰(�;+K?0���M_�O�B?4g�������W���0����p�a��`D8��/�jĂC��;����J�n�n��kHr��xۂ_���yb���c�]K7BBc��9RA���]�G���#Ӹ���D5��v�r�\�g�c��?��sL�V��� ��3�4!�pr��-�p�0b}}��A4��2�~��&�<�@Ȭ��x��HVȠ=#H�3���]��χ "5�L�R6���nx30�O�F��n�s�$��#\X�˗��e�x$�!S�E*�bݷШZ�J;8��~$����f���t���HZ�󁦌�t�/��?�:l��Ô4�#ۮ4�r�{I�uvu��1��[IFM�Y��ye��M7��?ى�汹v�>>x�<��f%�Ó�c��d�)u�NI�TFA|�z�J���C߅{��E��4(�+���Ijj��<3B5�aqDپ�๮�o����@����l��&7JC�S��5[y
��@?Ű��Ej���3|;*��齜g�Uee5�cR�r��V�9{P����Q)O����,��;KZ2��B '�Am���&n��gi%�idX�B=3��s���j���x���{B�{B#L��bU�Yx�<w���=U�^��D���N�����M���-䖬0�<5�Np���!}��T{)�-S`-�c�g!���9�;��4������K�x�@^2e��?>���}��R�８b�4@̈�k�8W6Z0�,�eS^��V�_�����N5�oajޗߋf7X�	�n��/���(*#a%�}5A����\��OW���B��FMF(n�x�����?B"'��~�b��cb����Q��I�r� 8$?'|�*����I/�@k?�µ�Фg������D@�ls>�y��`z��b�>>��}:�M�j��b�oS�����41���]�����o��Kb�Cf�+I������z�� b�g(Œ��W��}��8C~{9b\\��m���lݲ�{^��s�+��g_"�v.� +��.�\�O!l����%���|U�Pb��匕��3ឦ3c)�㠻��ݼ��|�RC�sU>j��w>����":܏I+>'�XV�6U@pL�zǤ2� �J���ƈ�*T�%L�t��9���+T8��ՙy�ʬ�f�r!6�E�KqӁA�	C[��%j{O�JQX�Y���I�O.��N�Ҋ�yg�����lE��S�#Ñi���LW��:�XMf���D�>F5�����[����ѫA��f�ҥ��T��J��/<�EI��76���ȳX*8���� �e�)��F��9�����A�=��a�aZ���Y�����_�59������_�h�Z�B�up���:&5^�jD�]ܱ�h�~f^�6zo�9f;;���S�*.ư��~�7qQ�е��r.�LF�e�����4��av!6rB�!��_�����>	�?4��iڙ���?���1�����t���6�7l�����%6�O��X�a덾�4��dhU౯ulw��u�4t���&cD�8
��b?B{�����#�	�,��Y�S������"��,�q�w��>J�K�`���b�J-S�J꺫C�Ԡ|C
,��~�?��{�,jx��ᑝi�,�>�?$����#�P(�X� `�\��AU��:B+P�-f���r$W���s�*�[M}�s��2H�L�^
�lZ]~b
���HW/U�`\w���� ��fwt�]9�W|���^�/U0���fOí�����ݔ{�Qb�2k�=w��P�O����[K>��@�Z�Y���Qh�*�r���C��-~�Y$d~}6��W�"q��j�mD�=�`�2�k��\��4.%|N�F�.�Ov�{N􆡬��,�h�8�6{l��R <ɑ����XOR�iz�^O:�B$�dg�7��{��C'<2��T����n�+�7$
����Z�?4@M�qE���1���E�RX�q_İД���s1//Y�gߙ�ߊ��Z��vI��ke��z�1�Q��!U��yKu���ԃ���-|���
��4�ȟ�y��@UNr�j�]��@��&Z~MA�-;�i:�_��K�Þ�3�Q�n���4�f���&n8ױ����4M7�~�MR@�.9����]gqh%�g�̳��݄�rV�?�f�T�M�e8�.�n�N�fg�G�����	l�M�������Y�h����DZͰ0�#g*�an�uB	!U�����r:����aaL�p���t�vaW"�6��_w��~����I�m��$�i��B�K�F1Fl��u�i�>��s^T��/��o�')[��~5������g�)�J���~l��U�V� �GMm<���k`sI���ٕ���*���R[H� �MӮ�tJ�Muiy����[��'����m\���<s��lI����6�;R��<��n^��>�-�4h�5�J�u�� /����~)7����H����n>���2[���|T��$P�ZL-�������4hڍ��moH�dcmg�#^��5�����DuL�~����1T�o�"�3×�l������Dk���FkO�6�7|��/�g� �k����a,s=h$n	���b�ᷙ�\��Y�J3)l�w,-��Db�,���r���=2S��'{Ol'���RA��O��֟�0Μ#A�L>v����3Lqg1�!�;��^N���WSQ�#�!��'
��C���4�!�����(Oj��ᠭ����c�n�࿅��>�o^��!�`�d!�',��4猊�ü��x��9�?Ld G�֐��O�œ{Y"î��wi�M�����=����'(!3��a��)�=��Vk����in���J8(*����l����O��eP�utt� x��+x������{	��pN�l�>��[�+�sD��ՎO�\D��U�{���*cz'����T|�%��pOM����;&�j��e(�˥^��ֹ�43�Oʰ��a�..y� �-�Ǯ=c�k,������pE�H�Kբ/�D��R��z��\Rf<�v��Rg�?5r�Uq��Q��N��|��kJ�J��~5ɝ;Jq��g-=M��s����S���~S���˾oΜ����/�OTkp̷Tӑ�Hl1�Ҿ8��{��A��Җm��)���♣�)?1�gg�x�L���ٝq�����$���/��@��|pJ�Y�O�f����gs����T�m�Ǽ�E^W:�ʅܵ�-Q�l��rUU.Nnlt�/ZZ�9T>����k�!�v'�$\Y���[�����Ɓ�׺wVuP��ʅ��7�N࿡�m|��h�4��d��U ���[�B��8�9���<�U�z�������6t҅̐�����ʦ�M)��}��Ȼ���X��
W�]	�k��
��/�8i�2�I#�6�%~�u�8Z�I�x��NF�[��7xS�ZHp�=��ɑQ�r!gh�i9�6�+Cf�O��/��E0s� ��g'l��/�C���"�sQ5��CaDYv<h�G~���W�y��P�Z ɪ�x�oF���8�E�@N��c��������oS��	�[��?K��� ��ه�Ug�=_ީ{|0�2s���uڎa_I�ll��b�gU�-��n���I0h��gާ�`��o�%�-��q��;
�I�����8�����_~�?�¤��Va��X����"	�7����'��n�a.�IP�A�9��#ʲ1��j�O���>��� O�T��Y�G��Lz�O�A���B�����՟��w�E�L��"Ot��_��5"p��?��Ν����N�s��٫�%H}��xA��&h���|��������k���G=�!��6i5GGwD���:�f�@	�%����"]P����|r��wk��B�l�G�3Y���Щ�>������}��v@��/`w��b�k9�����v[������^`r��!ەvGC�w'9O�pw��ʄ�E�jh�_r+}
t�L��vW�]�v3�Ѧ{���-_��}�_/֨���U8?�-��:�C`�Q�Wi��A����O�m��Z/W�
���Y�{�9�����q5�9�����6�0���ߓp���Gc�r�C�r�r�� �m5��C)Ϟ�ɋ��O�kf>�`ZP�W,�����ot�!9s�J,��@@�u�D��-�8�ehqI2���i��ncExB�L�j������`"p��'��SkY��	⟂�}��A}~S0Z~E�5Q0��7魩R�8-J6����m<����pYh'?��pu��X�ʡ�F[�ENxN�V�q��o��d���V4�=#��C�{%�@L�S�n��{��H�˻>\��|�}H�W~����0dI��կ�sB�/���4q*�q�3Q���dG����d�"}�ʁN"U���%$ps��6VZ�3�M� �hA`�}W��	��8����o~XFA� c�(Lb�iP�+zF��s��l������\�U��r��1���`�r7�4�.5Q�Hb�9~2��tZ��<���j��'o���Kb͠���(��� 5��(B��U\�L�y�y�+��"�egN�\ H͑9���y	���/dK���唉
��z�{[#9$�Vj������|ʵg~��/j{���Q�>;�H��Ȥ�{{�3B'���.�F0+=7���a96�_1�x����������{���je��N�D�K�r��*���B�o�j�j_�q4Da�?��3�݈�}�VQ |��&�~��T�6����@m�G>�:�>1{ڏ�g�V�8���Ŀ�%��UR�.������\mm��C�B���_cr�Yh�޼qY"U�I�RC�L������l�l�`&����&��7�֑ͣw�rzF��5�:�yܻ�8����lK�yj��VPj�����a�Դͤ���B���$��nG���c^��V���G�}8ea.�\�|v�ˋnǖ��A�LJ�s���llX��J�6y��۹Q��ڛ�)߁�w���tzЧ�澛֫�"&~��e/_|�m������JUQ��;\0Fڍč�V,�`��Rv� ߂}����������Ȱ��t��<k+����Sa{P��o��tHF�{�7!�I1���@��뉿dI��:3�c�(�հn�b�>P3��?P� ��g8���~g�����sb���	r�r�(Q<D���NUL����3��i�����4
��'�f���=F��ZlI�+�5��^g��,@�DQ�U��W�ߩ��>R��7w�N{�FT�?����<K�9*����"w�i�$����Z�%.�ފ�9\�)%0<5���1m0��m�bz���.�6'��hz�y����vc�t5�?�]MP��.Eq@����q�^l��s��MX�+���s�	Lˠ$�����/^f�����$
��2uW^��B�u�Ʒ���`���o���.�Qz֚���R��fx_�w��D@p3�9<6�c�P��ۣE��^�Å�M��5�.���Lн�TQ1� wG'V�W��D��nEt�6*�9��"�D�ˈz|�Q��\ڮ<�-����`���K�R�d`؁M���ؗc��&³�2)T�~���\�:F�1_S�t��4����1��l���*E��K(?X�����P�Ǹ�<(�W�<�&����- ��;�����	��+�9�0��7�/��W�E��J�̀]�d'���E�m�	2�� iNCw��c_�X��ŝ�R�(��*�1{�"�����\̋x�񅊔�0�6������>99�^����DAU.�0�NC��PQ�[����,����eZ�vƳ�3����W�o���Q�IήAV��D\�G�`QZ��½Ә��!����v}��H�wܾ7�e�� A�?�Hƛ7�]�#xW}��m5���鿓k��7�:�ucR�j
,��)��)O%���F��m�#�����~>��p�k��S&����W�&�{F������yv5�����<��J�/:��4
�w����@\9���~Nʕ�j��&4,�e� ��a�Y��0XgK������]��j�L�OX��QA���	�՘��[��LO�v�Q#�<}��  <���o��Ȑ��ߝdF��$���{VK�K>]�d��N���i����]~D*�bd$�'do+��#h�G��uH��d��1u�DV��OR؝ $x�|�`[g�ɟ��#�=�G9��X�������W��fQ�\����m=��`���S�(�[�^�)\v۠�<Z��ﵞk��50gpkD ������Z6�9�b��_��>�P ��-���	�?բ�$5�P�`wn �c�{����ވ���PGɷ��`d��޿W���v��fR��]w$�e�5 *�;z1ib@9 Ȁ�j$î�OT�i� O��ۋ�i�O�A��=�����i<2}�s�X-�)n�K�vr���С�U���A6ﳅMT吉�I�߫;�un�A��N:}�׏?0����݉��܀��c��F�QS�$Bˉu�m�*�~�V�͛��k�ar��F��z��=HRV��-���ݨ��[�t ��Ul��~9ѝ4!�W��MMA\S�҈�65�ڏp��`	$K_� �הq�G�F!��܅�lO'V�M7 IeO��XI1�Su� �A#|��;�A$�ߊ�o+���D�z��T�L쥬3��xd�tc���ّ�թ@�;���ܬЧ@]3��ؘH����IL3�P��Ȯɽ��(,��]����:�2)�%�����(��@nM\�d�,������@FK.�'�Q���|q���t���߃;�M^����%��w|� ���cS�`�c�b���gw�(�EWͥ[��:##8
��
�)TH
45;l+l�+��جW�zK��nH|lT�6�i�K��z�Ϧ��gT��~��M�b����}���Ԫ[U�~�;ao�ԋ5�k~ �L���1��ՃG�HL��� �I>Q;��ҕT������[�q�E��� �aKM+�w�\&���v��Q8�I`J��k��.붦&/��]��BYw�9ρ�3j�*��	�xޒO�4��k�7���]|d`��Z��7��`�I�z��I���T��RsI�N�^wttZ�Yk!��o�Ǒ��ҭ��G 7Rn��_	J��r)!�Vh;�0���~���u��O/!��]﫩�7�)��!�M�W��d(�j[�ITR����k������V	��0�֌�i�z�Z=@�Wı�x���?��Ş�W��_��>� ��AW�Cczk��Q �Y���fa5�<��bF�m�+�j6�Tg�p� =�w'L�}%z���d:�Ɋ�Ż�C����0B�s7�_I����{���5�.k�&�sg������$p:�tc�Y�-���֓����I�����|$[{�7���� �v�������g�`�	a�r����˧�w���G\4��0��S�
�~�J6w��[��	tZ��
�T���0O���~	�<O�3\�~{Q���	d\ �V��f
��
���CZ[(�?O�OTT�fˮ�b��0�E��"�긊S��;� X�R<�$n
f%��Y-�M��(u�ӓ֫�>�{��a�R��F_g<��e{l)ҙÿ �g��qO*�=\GR�8K���"Hg��gK�]0BnM�"��Sju
 a��6x��l��P��98��������i�=�6����:���
f	���\���,�n
u�R�4=@o�H7���|��9�_d���'Jn�'��dp�V�)�͓����j6��k!;���'u�.k��#�2}��:���Bn�h�ܐ�'^��`�xgM5	����Z���Ύ�~'2��H�<��AK��BO�j���t�Q�	C�5���pb}����t#�]L��ÓYg��_�)�����x�C,���G������"��A/��I������� 	�#��VI��)hM��J�	�p��)�a޲��-|�<|�
�Kr���~���5�	1�][(m������C Ɉ�?��'��" ��$;�縬^���=�K��@W�$�R�\ٽ�n�^�J�kw3���`Z[g�A3�6m��&��´Hd�ϣ�,μӕJco��Q�pQ"3�O:�	��@xUgG'f��$؄��9��!��O^ f��o.2F�=P�H�/���.Hټm�~G.8�)3��S��ጴ`��߀��>���7�9�\�>U�no��g�(������w��G��E���S�ɭ��ߋ�b&���X��@�#Ψ�%N�V;�Ǜ�@��d�,j�Q�>&+ 5�N�}h�����F�'i�����+���=&Q̉������u�EP�z�*ɕR�9��$�3`'� đ8�V���6���n�@�4����St�p��>jG~�86�ी:�0��)jGKu��7=,��˩D�bfzN'�U�I�s��v吝)H��ү��(t�9���� n,dױ�8���P������0Eズ�5�*��dH�PN8��VS�\�fWbZ�L>����)�8�-���[񰂷4����(h�G7��b��3`Y��z)�iP�ӓY �bI;���O�W��1�˯a�y7<5@���8Z�� 	R4�����k�������Ik��=�|�0^��gu��V^���,,�]1��^XԷ�CnVvf:��]p����~�����`oNठ����)P��NST`��~�MPw1v������ܒ�7ݍ��\�S�s_J�-BhE����̓�����4,Zcg���5|�^5�),�����J�M�"(Ū�NS�*�A��+�pb�i�f���������4����	S��^ �5&Z�,75S�W��ɗ�4|[t�� *��C��`��z�3�W�
\��w�tʕB:��%�n��]�,�J �b����l�.yęDfk@��e���Я��u��������j&�H�+a�@�����D�=W�@t��e� �IQǙI!��	�?p͋H6�7gv���ȒЖ��J��ϯ,�U��Z^������ 
����Z%���X���>)��*r H�������i���U։��(m���Mw-�Np�g#��՛���͐�rc���s;�Wˎ�f2�G9�;ϧ�O�&�`�;�1�j�h�S�oSk�J$������m,@t��l2��2~��
&\��	����c3����4p�����Z�� =�OrŲ^�vV����3V� P����0�eP0ͽ�St��U`����ă` gF}�4���i�	٢�Y�"���x�D����q��ĭu�$fG�<�CF�c��)�<0�O]x`�$�Vr�.�j����N�������I�����z��(C�Zj�+#k�#����_���� �Pz5kh�3�������9��X8�,�zFb��_��s�^�lԙ��(@:_wwUsG(pM�<{%X黪���W��r=�7{< �����#��k�k&R�x=5pvk�ߵ=���4jZ�7x��v���D�[��qOз�d�L�)�G>hx�J�e��	�✀���(.9�sբ^E���E�:8�����BB��h���n�Dv�I������S����l~�'��O�͞L	풔������`}�϶����~4�l��	�����ȽnS�Ep9����~iG���bgȕnHB�Gf�V� x;��m��h�p���,N�H��U��p�|F�ĭ�7[^x��p�w�	�}@�� ���ހ��P�ۊ��9d1nR�-O�pb����;x=qށ�/�GO5H������p-�tHТ�~�d�}=!�_��-K��H�=Mޟ�N���5�����>�N}�|gP�'A�"��b·/S*���ӧ �#HA�(�c�
���L���U��R���.)��m��m.quل�m�I���zt��1K�)�c�N��4��k�⿞��Q�z��c�H����2��yX�j�Hχ�=���̤a;�X�uY!O3(��e1N���3�$*-=��W��]J�# �1�����W�ε�XiT��t���2Wt�2�FD�*�e5����F����@��v�KC�+A�ļ����/��*�D�c� ��]P��u��������&+!�����:9��s1 M	�J8��H�[�����������1[��a�۫l@M��%�񙲍P��6q�k�+��C��M��YBMY�9�jM��Cs��,�fDR�u�e��>�[�V����it���ePE���6��^X_߱���V.��@����҇�V��S x�&tC�F�����aZ�8���T���]�nc���Xd��r˻��������U�4���`&��)W0���/��T�T;�^s�����3�A���#�R�l)�bp��|��Q���	ݘ�� �T�)K���<]�vg��H��o[��k����
���X�%y�G��W1�y��3E���"�әpo9V��og2(4f>x������ǫ6���O]>R�5e�K{ff�tN�L�t�iwimv����^���=�'�6W��&'+�D�-;뢢��
�:��	���y3ߪ9�R�d��d��Y^�H)��������瀋u��â��Eƈ����ϙ�[��5RN���p?
L+\�nx��'���R�ߒ7ݳ]�xx�P��(����~��1�8�2�v��m�&��/�H�D�J�N�]P�d1�0�-1��k�P�a�=��Ҡ����BX���u�$3.Ss� ��b����Τ�فI�I�1���
��Ơw�N�㰷���r��T$+�@��y�w7W�5s�\�Q0/}ƩR��Ƚ����)͈�[K\�ƖeBnA���$6i/�?ϰ��).�u�L�rj8�p�죡H�o�a����������'T�*-�hV+�I5(�"S��B#�'Ĵ~"��J��q��m�o1�!TJ�x���t?b��6�h��-���\����K��S�9zuz����jbEFE���3���Y�4K6�������3K�1�2�̴RwP1�-��P� �{�����������T^-t���$�Y�Gv�R�d�y��e�Ԋ둖�e��ZpM NS�9�T�8s�r�Մ�a�9f�W���+S[e��ۘ���"U`i�b�\J�Xz�[�;߽�7���6�{�#��a��j�Uz17���O�z�5���>� iĨ�1��p2ݥɊ�D%��J8~�����)��.�����
b�U�_@���c��-������.,���� �F�~.�|���~6�$9�M�|�>��]��a��~���4�6�ߍ�lS|@	�y^ON"@���(��=���o��WhRMbrm@KCl�0���SҎ>�Ft;�r׋��y���P�>�}2�x~���!��|	����OmkT�O�&_�g�c�:;���)��O��h=\N�ÿG�O�V�n��ݰZ
���l�Z��8��(5X�8��,�E���C�bK�%=��HK�Jk��Wxo
]C��A/h���bz�h����b��*�/ۡ4Ե��r9�٠�Tt1����Q����N�Ɖ`��^�rMz��<r�b[b�Z-�ns�E�Q��O�����#�=�1�+b���"񚠠 �{ �VM9�J���"��Яw/��̄�j!p�W_��c_$Æ�Ћ2���n�R⪪jG;�8����{��W���#�{��娑@��?�;�~ LUE'{m��̓��	�`�+��hѻ^qd<���0�
h�v_��Z��Ҝ�b����$72��}H[K��'��;{}"�K��M[��S��=��9�{S��(dJ�6Ub���*6��e���J��[!
�<n�b��.�Kw\ƾܛ�޾ݷL�H����f��s1pi�&p4ר�-�?61����z�7���6.��e��>��r.D�?c��d����@�I�w�0"�-,�5RY){)�����_��)��a�b�ݷ�Y��m�w�29
` (�F��4��ȿ�8��p�eha�)9���X=`�̵x�Ba��, ���FI'�m4���Jr^�i
����n�j�]k�F8�ۦ��mh�����zr��s��50�31���Fz��t�����L�Ϩ�>�C�
s#ai�f���us��yo�G]z�͊�JJB��e/{n��*�}H.�n���H���v6%k1��t�X�9����-����Ø8(i���@};��������P
���N�Q3,\� 6�N.�O���4�ݽ1�����m��hGBx�,�@��4|[u|0��'�S�?e���Oef_�-|ҒX��>8JO DmX��PN��ޚ�,k�녜5+Q�3��-*
������`Mw�q����D��	V�̓'\n��̠;���-32p�jq�7��(���1ȉ�#-�'\�8���g���~���A2Ƨ����j�*}5&e�!�P=�C��������̝���fϦ-K����|y�V�,���GNv.����Xٓ�5�����ҽ���H�@6�(�Ra��]syugW�LJ���L�ƦШ���9t*�9��b)��В2�TOm��~����z7���z���A�5�J��^I��M�><���ԓ�p��;-���(�ۈ,��4�42�U;]�q-�����X��s�ʄ�{|�˹�"��v/UP�K�e��=�Ѝ�\��E�}���x�k�t�Ec��U~�t�����彘���Zf P*N�� �&�\�!(R���	��Ef��=;�����Y�ߒ�-��ۓm�x_�'�[m�0��1�:��h��@�z���6���|���r����RI\�N w3T��@�~Z���l����!.�O�}�v��E����%�� w��P�����y1����;0yƂ�"��(�C���8�7?��k"7ҵ|���KP
��#����4�QV�sv5 �	�b�pҶ�����k11qH5\�_�*�:�
ױ��Uq����G��)Ե �� 0n�܌F�6gr�]�r[���IbE������U��itsZfw�l��<F�7��ঀ�A��I(/�r�����Yrv�����(����7����4V����P �n* �$ ft�-Ѹ���<�NâeK�_����$6��䵓;P�ê�M�K`ث ��T��C��םp/::�/�������NBJ�%r_�	X0�(�ŕ&�j�fhXh��� ���c\շ9��Fr#D���}_,�2����n�Ի>����.���d�� ('�����7Àp+80�W�5:i�K�ʝ�_t��~=Hc��p��>o}�!#��Z�, Jl��� G�ܓ#o���1�Xס�'�Øp�����s�QU��c�$��i���?72�o��8���2���Y�:4����`�Uˈ���������1A��԰-�x�w�f���e�X_����)S��$�-�ؾ?yO䒅�ôP��Y�'�J^ѻ"` �(�/﷌ơޭ��f��Z�,U
�vT���[^��0u'�j������JS�F������9_��tϮ��\tټ@Ѽҋ�M�IB�ˮ�d��%�K�2�R����iur��p�+�������A]��)��+�[p7&�}�;��X31��B�i�w�� r�5�d^w�n�)�G��&a�����9�G����[�d�(i#�u$���/�p?�\�yiϭ4%��*�Q��F6Χ���󣏢]�CtT"����ӵ�66�� "���e��rv�t�;pƌ�x{��Uz$Y��s,�a]S�d¼Th����?5&����
z�3��� �T�?�� ��@��#nJ|-�#E��s��i��N�)��Ĳ��U��`	-��-ւD9`��Aт�wB�6];���R�����,:��!��kn��R[
������?qauYU5�&�E�!��+݉�&=�I㍷�;V]����;�}�iǚ/2�o8�n��� �-���z����=�Jeuk��ZT��s�F�m����/F�P�Hk�qA�� e���W9�^3��7R5o�$A��ʙ����v�b�*��0�}6��}��6/l?\?���l�᎝����A�ɳ��n0e7�7\V�m�z�E �y��t�J�$ٹ����\���`�"�}Q���[�~����p�:ⴟ9+��4������o�,� �ftP�1�g���n�Y�?�9[�j����r�z)B��h�F�pYM�U�����9So#	�����Z!�^�q�-h2|��eN8�|�c.���?�=Hìu��R�	�������%+z=!��V�����SY��لNϸf@�r-�Pq�}w X#��"/-�§��H����^�,EO����3�\;�,�l�[�a=liD��d���!���zjo��B������т���՜�=bg	:y�B)��-F�*��}U!,8xM�c@�G6�Ƀ�w�?;�V0�S��ʪ{�W���>s��R�����!�y6)��%$E�� �ߊ���(Ra%��n�Wv�B���yz\׮h�;%���l� PT=�L*Er#���pI7&�#�wӬN��	���� q�K�NPO]w�X$���Nl�.�|���z5k@S�7�0����eN�x��M@��䬱M��Stog�N���}���kO:g��^`�F�D�&��˂Ǐ�o-���J��C��#vA3D�;�W ��lP��t�`l�&�ߗ��x�n�$���0��G�G8aPE� ��	�P�R2��a��݈�|5-�o�PV�?�jYl�"�gb�sLI�4/G���Iu7l�lM�ڃ�z�d��/�g�Ŝ1��20�yz0]=r��A�b��~u ��� 6���бF��Cr�R�]t��NF��~K����˥��1��Р/+�m��7�!j#}���#����Q�4H�>�+(]�d.�A�+�,
 6�t��m@z��S#��5�L{��Ƚ�+w5	��~�Oa=r��X�	mҷ�K�����5��BB	@�%�g_�-i�w�2 >�[�nC7��\�qi��&_[c?!�/A�~�4[��������]�8"o�D�Ec>��ӠV�񇞿�n?���-6O�>�=
�{ǡi,��-����� ��=S���1B�!��ǆd�NM���WGB]�֔�ҋ�K���df8)��h���iPj���'q�x�m���o��R��?�V�48� ���)�>�Oӓq�~PN��<�2[��Y?��də�erKJ!ś(�,}��q��g�72;�9��<g{�Q��9M��+�ө��t�W�i�V�s��AIܨ�\����N�emX�tɯ�k�����Jn]P�����I"OC���g�u�O�ۛ��\:����PL9M��ʅ���>�{���Ț�z���X�{=c@���n��5b�\�	���&��M��ؖ:J�R�Y�.�b(�4���Q���"&|����~ʿ���8�))��,�P��9@�%�C~��[{&\i�%�mW�	�%z��y�^+�:�P�b�PP{��~��k��Ж�(3ZOVڠm 6E��ƶ0Mn{�ߐ�U�*�q'�P�b~6@a^��Jo��C-}����w�e�6��-Ux{�y����l��M8���������#�<s�,RT`%g�V�/�3����~��V>v��8�gP�(B�т��A�$������tZ�U�<\������p���bw�`��iX����� d
�bƷ���Iw�J�����<i�a�F{)�ݻQ��9�#"�@KF�U#��uꞩz<�b�0� X�~��C�Ld�P�X��4XĜ��n��a���M�t�)ֵ��LFX�4[
��A�Cm@q�����S�VP�#=�[2��3{T�!�����kroy�WN��I-�'��A�����N���J�����-�%�s���!��4�ŹY|��:n�L6���?��^��HM�&!c���R�V������LM͓QK+��.e����>VKn����Dw��'���Y2��A��Gbz�*ҿ��)��Cl��3���Ra����u���P�HX����e�@�}�;l?~JR����텈X�!�	��c�<�={���)�/�3*�d[�E�qP�A$IV�MlP�YB%(��$�d� ���@rlr� ��᫷	:s��q�����̑�ߪ����޵�:I�&���U��K�]#S�ڲ�v&�^�W�[�W�ڛ��@b-����o`-:���R��^51��G��^l��F��ŔJ"��S��6L�K4�,5�|�hkgRe���LM�of�Md׿�T�V8a;̹P�+��r���HC9(����VV�Ȫ;� tb�P}����@6"ⲝ�ۮbU�v�=z�����	��G^��$���(���z�夆_4JVu�uT�I$�mdA��W��>�^�	��<L��r���['��	�)�>:����`uǊ�n�BF��N�S-!06�Vm嶐�.�V��yy^i|;��lS ���-j��Ĕ�cY��]
ȣC�����o��7�l�D�G^�q/�]U�{�=��(=4��]fC� �C����Ei:I�Ƞˈ�N�ƶBA�r���J�V�U1�:�D�U����(W�e����M�1��I,Sq�|(��_,��c�ҩ��W�꺛@[?7���/fu����T|zI��\c]�O��.�f���Yk���./ۺ{���Y?%��y�:���Z�t���]stqY�rWI���5��[�t�i�-�%��7����0?<�{d1hWW8�V� *����T��Z*�j��,��`���&G]F�+�|�J��ߤ�����F���S�
#��u��5�\[�tm����x�A�^24�ʟ��r�`@�b=�![�6��)����#{��as𝕤���lm�P�hR�����C�O�&`�}��D��W�Y_I��$��L��m]&z�>�1L�f@�ٞ-&�i�	oꏯ\�v���o۝�q�4`�.�t
����P����J=�l��T��N��]�5�.uʦ��@s>���v�
*RԄ�IAg@E2��� D[\q�(�x+�^��p�d�(j���� 4��|�U<�K�F�ToLn�������9c�ی����3ܪ�N��9�	�&�Ft�90`u�a�U��ЯuS[�$�T�p��|\2;  �z���p0�T[�uh�,�t�UƠ{a��s8g�eu�LH"PO6���\��hӶ���6��\T6z���v[o~���Z�\����L�n��]�"@��-6��A����=��!��Ƿ�^հHK�X��!$�!p�{K�s�V��Cݟ=��a=�)�ҽ!O��,�us�4�@��A�;�s#���~S��إ���5�ߏ���5I_���*��JO��]rm���p�|�s�K�g��UmV�B/���#=#p��-�fн3�%�.[����ڢr�rΧ��]��Ռ�`=�MAj�����n�0�����uӕ�v��zغ�ܬ���HA��.xǗ|�(�8�B"*�?���j��	ڧMl�D����PS�?m��CM���m�\.��q߁j8�r�	E��Q�P��j��3�+�[@Y �o(�����ss�h�6�x��0��@���E��H�5���B�r�����W�����3��GG�:��u�ſ��^�61q�9Ά�v6�'�*���Ҥc��B�2��L֎���P�0`Ư%V�T7��Ջ��2iVC���d�kR����#��"�q��izm;W��=xS3�۪S���G��{Vo��_�ze(KY������ �V��Ƥm.T�r��i7k���תV|��O���{R���\�@�8��R&���EA{ �.�,�F&�W�-��=��V����*�����+6qn<9?���~����c���Ʒ� �G�G�EA
��
(�ʊ���*'��M&;YFz��?�nˡ?�}�_�Ư)Rw���G�MA�-�(K�Bo���N��_��/^}MX-���/&�_����`�!8"�j�U��Gɒ��
.º�3a�\����� {�ڏ�������kP�/`;9G��sm�h?J-Z�Y(C�z*�ԣ�
]�=4x����A�����	�215ge���H-��\�9�[�jO-?�JzX>>捖���s�w̻e8����{��S�?D�C>=2�唯/�:����A_DS�M ��eF���2쬠eL��a�����]xc-���Xdm��lrQ�4�T�J�#H��.3�Qrd��o�\�ƥ���Z�"}��~�\�o��ԾY�bD��V�����]}�B��+v�ЃM�c���Ք����@����S��Z1�&A:�9�~T@�Yu��� �P6|��+�o�K��VRR�pUO׍���ݱ^#���s�_��Z
��Mr6�^6��~Ovv�͇�����O��֚4?1Bʽ���+5U�̏�����(`j�Z��9Z^2��D�<Ӟ!X��j��,/L����W��n?������"'s��oQ��T�E���Y���v��yR�a/ s�_��3-�?5���5$��+yV$+ą�|�.�
��5g�}R���O@ ��5@������%rv-�N�d��r��+':@[�̿�o$��I��ICs}L-�^L�;E+k�j�{L��z����f�as!����r�
,�RZ��uT�f��
[_�Il)P�I���y�B�H5Au4� s�>�@�K���"~wߓ�c���>�� OM�)�`�Ϯ-�Y9
�[!����aK&К�� �8� ��G�	9O��&4ƾL�JfD�W��J��5���ڈI.�~{v�MQG1��:�@�]/�Tuw&�#w9�)����l]��>�e�Bp�4e���[ox�r��r��톿�r��h����h�
���A�p�d�T�S9
���ߓ��U��� <�@��K�P�� �tq�p�!Mx�W`���K�x���+$JtSv��p�21�AwQ����7''�`���s-�4ȐӞ���N_	k����7�(|����*Nk��J/Ϸ��Q�W=:�]�����o�`�E����w���_���|�����sE�/�)x��KR_�⤎�M�([��@��΁����Pz�7�e|x��;�[����`�g8��^��j�#^e�v���7�$��R�K���\V2agC�<���G�4;D�����f�`��]V��:qXwgV5T�\�55��i��`t��F����`���������ﾎ��*9 �4V���N���^w��wrT����rK�~K���;]w��~]���I2�dϙU���Y��ȿ}����F3C3�����w�t�w{Nk��UV?G�妻e��d�X?��aς�*"�i�;jWo��
�I�P��I./M*�3PUefF)H�{�2�TT���]�'\1w���1���㇏_��RP~T������Jz��#�P����O7{�Qr{pm���7�X>�����wd�!�Sw��k:AbySS{�o���ћR^�H(����~����c�:�j-�E��,�p���r��ͯ�z�t���4��l�}��\Y�h<�� ZƉ�L��k�N!E)�l�K��I������?�z�7W�9>X����)�_-G6�hw�sf�j]�nɳ1�KT�З��~=P����ޛv�Y�3�,��,�&��Z��?��	%�i�}C��ۖw�	�̈<{ػJ�Z@��g��8�?_�[��1�avCL#z�,[B�U�G��4�^�|�h�鸋���C]��'��5�
hn�[������yt��Z�H�]>X�q�%V��p�9�T�(=�*��[��o���%�r9@k*Dt}5���f��[��7l���k:���Vd�^��aƐ��Ly���e���A�ٞ�e4����O�}��3��ϖ��M_B�gݠ�e��ry�r�c������l�o6�ׄ�UG��2F�� P��9�I�=[�'q[^�9N��}Ϩ����
e7ڛ�&F�,��Λ�	�<��;魪�ޢ պ[rq��+Z3籏�V���@=�&�mλ"��Y�D�<�����+�cfU	]�ː�Z��7[ �\o�d�׌gs!QG|碟z
�z��J���R�\���ZQ���@?�2�����23�9~Z�7��D�5Q+o�;���.��|#0��dϏ�)���k�58�}Lh�7�a��^�+�7X��	��}��*̘���%E{j��w����1�j���9V�~ӽ���A!V=IE2\+:���i��L躹��5�=��N1�:\����~$��x��K��Uf�]���+���~�k��"咱�34����Ɨk�����$��L ��U%�Tvf:q~!S�⺦s�B(X�:�nU�ܻ���%��]TܝbD|ۦ��&�E���&�墁�E3Ul�&���p"�78�: �^���VQ|�\`���O�Av���6*5t�O��1EBߥS^q�z�~���K}2|x�s!|�	��n�-��rwɏv�ʎޛ���<��\!�b���$FH|�@���s�Q�dαq��e�r�`��N�s>N�
�����l��^��ް* !���6nzM�>G�Y��{꘵�:��2�����^t�9y5���8����)�"�=د�O��@����S�����	/�:��^`�*�Nxb��ː�T�hَw���I���� ,X������ 3��.�l�ɟN�мe���[� !!����>:��4Ej2��j�px��� ���rq�rͤ�`I�����\{�-�n�E#�'�o����EύJ5`(�������)�[Ɯ7²|�������#��W�$�:���3z�D��ݡ%�!Ku�w)�w~�}]���9s�ʯ#D-�
��X?q`GC�7*+q>�B)�n�����$���$�sbLh�P �� s�Q�7�%�,�6�vV_|��6�w>O�o����a�3��.��!5֦��o'stp@��$�q�S:���!��p����t]�@��d�ޫ� ��H�7[���0CA��9�N�D��6����akL�jq�?���t68�tb&�7��W���m<}�'�����P�cB{F�Et_�c�>��u,p_���|�S=�[��sb\Z���c����7`Dsi����;\�s��i��:����Q,^�%D�eEWYi:6hhZ_Q�֘�G�:j����&E�Ġ��a�ŋ�/ro��s基V)�t	E��!�)O��M�\���p�:���	Fו���'
�x�@p�1x�*A�+�I��c$Y�#0�͟ݒ�����{�٭k �4����x�d�Yq�4���$q��pn�O�R.�oU�06["�.7�H�*��}�4��T?TCT�F]tx��5'\�:D^���)�0�H��/96�**�����3���s��Y�,9I�����G�!�̈́JWz�Q�H����>�
�TS��bp4@ Z�k!�����U-:�ne����,���1��$�؀�p��d"𦏴�L�[T���k��T�i����z@?����~��{�^��p;7�t��H;+�D�������l�[�(X�l��8���]ÂC��gA�@�3�Ȕ��\�s���=��G��7v�*`	vy�
��
)/��U�R�Du��͖j�Ư����z���	ae�hx��^"^]�f[���}�o��H�&����W�r���?c� ��qr<�h���zt����݅��*���L�g����^���y���7��b�ҵ�1� �p��/��A���W��]����Y��R�;��{*@e>Ȉ���}
b��F#����*�>.w��:��7�_�?ގ팡�Bl6�]�]�_�*x3.|qgX.^�Cx�򌁴��!"������}��}hP� �m�˯�Z:��r Q��~�ݭw=:j��#�o�g��[YFw�b?Z�R�g��{��j�!v��=�7�����&��}�{�1p�E8���6n*�i�y[��-������r©d���m�Kˏ;z�����A$	nA^���ū���M\#������pNQ��C:�}�~<� BC2�VUpfy�U���YwR�rH%uMٮ����48��z	��H�׈wB���,ť4q�9�T���A�}�s����l�_�'���q$����U�Y��"��Qf�v�ZT������nF�Wg�6�ƶ�<"�	�>HB�NMl��S'�ϗ�	fqX�Lޱ������x�c|�w#ls-'�mc��G隿��ʺ��%"g^SL�ߴ���6"=���]Ϲ���s�3�f5@����^x'�^!x���)��<T+���i~�j}�i^���';]� �w)K'�H���F��i�1��R����"+H�p��]yxK�%Vg����f^u+��N6�2�e�?d�tR �Z��4lVk��J�[ƝG|�>��Í�
�4tDmN����F@����ߍ��Ձ"���A����R���[ < �U{�L;K�«�:=�����+��xʼ��S^4m/ZiCٙ�F*Ȑ4��J�<�Sy��-�q����g�*j�?�����|�y��.�|�A�0�ZeS�33�QQ�F�=���<�����s+�g�/�ޗ��s�s��~_.)9E���Å��N��sz��5�H��j����	�;N���KY��C�(�)�:�:>xc�ص�0^����s�b��<%�_;0���"���-tr�|n�W��+�7~�$q50�mu�'9��x\<���
�\%|k�氅L˫�؁f�M�-G��o<x����l��k�}���Mk� �&�ή����-��G��Λ!�sp�d����O��]됁P��TMT��9=K�n�)�{Z�6D?SС7��+h˳�bdg�K*,�T�>3ثg�k�[�֔��o�c%b)�g���f���T��8�u��+NSe�0��e�=�����x�5cl���(��r�2~'�Q"h�A�sg��@Ǖq�hs���㲶���Z�L3�o-ֺ�=�ͮlr�ݗrf���C�ٗ�\a{z�"��h��G�������^%��݊�i�G�;'[����ζW���2]� ��r�L�A7z��=����deA��	��@���DX�E�5~)�&����R��u�+?-6MG�E���W�-���x�C�T
�TȦ��SҮSf��|��eTH�c���])��$Z�> J�Z~<��w�n~��.,��Lc&`	�#�˾j<$X�k78GI6jF����n��D�<*��!��wv}�$��)m�����m��Mc�&:�$7=�Et-�b�1=<�y�o�o���Uƺ&�V/����!�Yo��^���p�o�AYb���"��u�U��d�;B�J@F����B�㍬J�F����qȕ*����� ��:@��.拎hѓi	��� ��}�_/�l:����/���;����@N����*���߹��kEL��W��zdɍ����L"ާ��I��> �Q6,r���<�N�ކ���֘4�j6|��ljW�R�.�d#+�WJ�e�_��L9��nq���REG�y�x���AT�K������;޿*Y5s
*zL:45��d��R~���E��º>�SCY�<p�%���k>P^z��
.a�S�R��J��; ��xF��&_�@9E�����2�~�%�P�k�K�W-E��|�Q����Pd>HT��Pv�9��g��T���m4N�QQ.WL-�M.k0�g=��XCk2�>c)L0� ��_.�Dl�p�`OL��� ��-��Q���[�p������17%d?�fd⿪�:��U�ye�`ğ���P��i5UU�[JT�I/J���¥Cz�h=���ߕw��n�ƎM* i�؀`�"uL��-�-U�cl1�x��R@��-����c�@f%I�u����W���Ų����晞��p�^}��o�1���ͲT_}e�#�ܨq�Y���^9�b�3fŁ�,���q��X��)�@���B��Z֕�aѐ�F���O�k��(���XX>�Z��ڤV}Iʲ�𙆊��{U�{��k=��,�7�/ ��I�����g� ���A�VA"G����agd�λ�P~��4{����:j7�`,����|P��k(�;�T � ��� �Af5�cWF�Aw4�|;�n�e�֟��}�4�h����������ye)9Ջ>dl1�B����5�8����3��*?�����x�c�-ݼu�d������M�J��E�̷K�:��یRK�z�6J�Z><w�<<���o�W����[�fu�E��u�z��!����p���a�뒡eͩg�1r3y���Ke���W��$�/�rQ��q.�nt�>�H��e�p���H���d��n�0_Wֳ�!!���ff��7d��T��T�!ƿZ6��uv��ު"�[����l�c��r��[��r�n�j2r���Ϥ�@,K$��v4�{�0r�X^&Ř�7��	�|�s���˜��ʪAu,��m�&f�-���۶��� ���S�m��Y�܅.�#E�y��>�Z�^��M��(-��6G��Ƹ�')W�/Z:�, ��)��/\Ю _���u�D��OsƎr�T�q1�c�73߄�g�2/��<�����,޼mT������RafU|ck%Qt�B��������Y��5?C�W\Z�;�w
im�;��W���������6���W�>3L꡿H�-��{KɃ���$���5X�F`q<~�yË��c�����k��� VY9��h��sn^���7 طDv�7���FG���n�D�i8��o���TR�O��M��w��^��w~n��! s��Q	������F�I>\�?��ɦ^���%��k��	 w�8�־s���^��7c�����CJ�.��r��5�L��3���O[�>�26���Ƙ~�O �<S�I8�l�`'�y=X���Ҫ�{G��Z�~~�m
Q�t#��0��Vڢ�?�/�9�̈�oKi�,�p���b�$��N��	�T	���,�yw�i�kH�J��թ��s0���5�w���~��WK�(�'GZ��#�"〰�d��l�y_�Y6+C�'�̫E5��4�|�>Ce����fcC �������P���M*_�_$r"z����X��}�����i.y��N|���X;ȀL��7"�DwVM��Q^�AN*j��̭��ʓ��e�jqH�m�֝"I���Ow%��O��� �8���s�����Y"�������fUh��-<-!!:C��!:W8���Z�����6��W�?�;���2���H��/w�&�0�B���`*
Ť�-�:�����_�KFJ�/�8UC	siy�P�i�.��^�훖�/_�����0H�A�/"��	��lǱ$�B�4�nw�дn�c�m��-D�x��I�n�h*���{�x�<<7���:v��mk��^Mld�E�	��Ye��ɧ���X����}r[ꈗ8�RTˑ��E]R.Z�M1۟�4�S�C|�$C�µ$;tR�c6Q�	
��@�MFj�v��+��>��e�4�����o�&�k{�/f$�����R��~��	�K�[X���i�<jH�!q��N���7�:���W$�g-�1��<7'�x����*����R�Ɩ�v7��!���nV��`[/I�c:f%��VW�%a(m�Z�8�#l)���b�Eb(W��л�~AbjE�D�"/�1���.���N�\��}�#)�ϭ�����������V}.��?�+�ۡa餸���S֤��ڦ�b(k^�[����f���S��4����,�	=�o��yϋ�}�q=���ݷh5>U^켌Y��]����c:ж..��@c陋P}"GVk[e�i!&�6_�_1	M`g1���
�6��Y���M �Y��{�� �c���F��.I�F&V�	��)@��$�̎��d_�ϔ�%Kq��]l�n#�L��(j�m}:~P��������T���T�5��`s,�X[�<o��ݹ�Ͷ��90y3l�k7��/W�Q��0>�S��T��#�&���D.8BUo�����~�q�_Nl��r�K��Qtuv�i�4�1Xm@�� ��0�k�gP��O�8�4spM�� �r�։<����Cm%S-�a��{�|�	��OX�v���{բ���Wf�t�A�9q���r1���'���\r�EO�T��TCf����D�{YC��hRz�tLFw��n��S+�<5V)���4� X�6W��*����W��B�z�T*4��|h�BO�Ke����"3�w�
���m��?k�^�$8 �N1�U0�/�c+�,|��c�O��ý�����"ٯsQ�|e�ËD2�7m�*��*J��&s�Mwźљ�vTȲ�����޳J �߀����hH:���ټi�aP^�B�l�F���9��&톾㶂����	��9�Z��ml�뭶�|���0gk���Ƶ7(�E��h1��娯H��mq�g+F���)�Ⱥa>{��L�`*9�k\-���q[z�@��%t?��}�KRoN��\���#a�r�\��p0�F�`��H��绸����t/�>�%�^�I}�� �S��7�����q~�¶b�"��,���~�:2 �k����w��L�&�6�>r�(���,I&��Ȓ��M�A#���(~W*�V���R�WITE�0 ����$�5�J���6r�Ep�n��%�b���t��P���60��qa4�s+��U��A!���]��r�,�=
��8���Ơ�vo3a��6ez���� h�(�P�em��8�<���Uޟ�%ǆ��M?�u���w=�2C��f�|�>����%
gJ�{v��� ��v����C'�6�Z7+/����
�X9�D��u�w�^���l��f/��B6���)�Nkl9������Y:�ΙK.=|%b�RD��p1��ﶬt(a�S���\�iHK��ĖZ���{���i��DFy�]mC��(��Q�� �!c	K'ξ}v�/���]�X��aC�tE�����+���4� K� �F��0 ���p��O����))"2�N7l�0oϕE5��w�d+�R��16�aK鳘f
Y f4�AEA	��]2�	Чp��V�'�)�Jʡ��Q����^�(?�>+�2��_�;�a����\|���.�k�4���\M�dbr{<O�7��P���k�L���]�zc�e/�8��Z
&go�7H�`��B�t�B;ػg�@������i#5��J��^ ����b��B�U�ّ���u傱i�C~3���z��
9�;���?���
�v�_�6�>oQ.zK.��k5M��i(�߄����7z	��������	/�k�w��8<f��c�+ e�\�m��)+l<�̏*�g�40T��.* 1'B�m+ ���W���>3X
Ҷ_H't��Y5�G�����>ٟ�����+����ၾvr����Ĥ�9�A��O�v�v��po�Z䧍U^')�O|@���Its>ޝ��\N��� 1S�|+�i03�T��\������LI�f��KVf�K��K��]a0!�C�bd���!pb��p���lȁEȲ]�/ѡ��(f�)T��L��y��M��nQ[�.�� �o�B�C��Aw���0RQUU��	PO�W�gj�n� 92��#�~?M�O�$OY�|��
f��:s0��C�x�b��mnQ *A���p����P��Z_������TЋ��j�[:L|�⏒�F�QQ�Y7���>>�/���!�_���hhv������oWu��k_�L�jrZqڴk�9�\�2T�+�.�v��jG��h|M*���Md1��v��9�[�x)��B��u�td6��� �����|�s>���n�C�V6�����5,�O��q+�Lg;���K����³�n�۲W�9����hv^b�ųڍ��͡>���@�F��D�������[�[d��[��mh��憦�/S��ͩ�����23x�{�D��k3��H��\��|+�6���Ý۶x��~��wC�B��d��q?G��������Ӌ���\,����x½������Pu��l��o���T?����ٍHC;*����t��[��� �O��f��r6�(��Qf7�oN��v�s���U?H���[�[>++?-$�8f{����B1�B��0.١bJ��xF�s��}��tá����|�C�o�:/��������J2�6d��΂��ꆱ��֞;���Q^q�gdq�箋}��@�r(�oS��\<�`����Z��(�Y��-u������B� 1����0��S�o�M��,jU��:����#�jV�%��YL��ߕ�R��)��ۦ���֜�M[[�QJK�*�yֽ����?1 �4�ϧ��z2A_�pP��ɩ�i#q�`M��7o�+w�_��Ov֩w,(�o���}�v�mS^Yy�Ff�G
p����0G���Ƞl{�3=9�Л�y�r�i5XyB�j�y1-�w�ך�w�-��&�]J��o�-�wN�~�<E8�ᶍg�`4�?<Kk�c ��J���>t�9/�afo�.��أ-7D�l��H}#[�T$mb@�Jʔ�z������\L�k"�Qc~�m_�/ᙧ������$\'z���Mrx냄?��<! ���\LvߘC�v q�v`���ȩ�z⩲l�ޤ��'�>��q����u?u��p��@cæS@��ޭ{�@|}�",%%͞���8�;	o��7	ݡ5�R��6��p=,4��A����z��:���v��nۿ�X9\U6q֣�P����C��-������x��莴\rۃ<��?��>�G��~Ҙ����h5@��H05#dwuNد�6`�T5�_�}�ۧr]�h��\��S�K�6+�(��-��_0^q�Gm�".����g���7��z ?���(�G��eU���4�#�]{U������t���m�_���¯6DE*���,.�j>=P�NH���	�_�����K�����t
w����穼E��1ވ ���̷�:Ρq50�w4�;��qISb���E�j�#ߴ��ڣ�����׆��ARf֐\w�jm�+�����Cɿ��WWS�h�1nq)�<2�hop�ֻn��CzB��P.f�Y���5�:fx����|�%�Hǘ��Ø� �5�[<O��><�;j���M8A)B���p7���k����H�a��)��6�_�j7�~����EG���~�E�m��Uw�~��x���1b驨�b(�#��#M�_e7�����c�& ��[ڎ�4��]X퉩&���󿒹ZӐ��\B�a"�X��.���_#|��f,� ��H����D9�V=�ت�7IqӞ�x����F��}��Lj'�M�繯/��K	�
ܡ�?- �z(�i�e��V�1�D�+�꺉�A��vJ;o�X�9�Y�)�9��P����KB��+�Q7�vS>��#�z�\�n����^X��cl�32��>:l��<?��C�iG6g���\"� ����=S&p��/�BsM�50��΂����(o� �/-����Y9���DFG�����t�ܐ�j��ZU\Im�[�O?\9R�ȑ%�3���g�HR�9�F�裩�n2�����Q�و#�� c�j����YFؐܯ�s��I�4L�
�d ����|$~��=qd���ڵ�j�_:�0�1�����E����#��˛aƤ�#t�27L;�R�۸]s�u<��im
:@�	s8,Z�e�<R���_��'��p��2�����9��G���OVE�����?��J������v:���`ek�;4���r�H��w����u���~@�V�CAE=��ܞ����߻G�;)�=OO�?�$ ���Uj�]J�����UD��޳(�s�U���2��_B-qq�{��e�n{{b�1���YV��yy�&���G����?�
�ߎ�|#ؚ�U��(�G��h�R��9M$ BBtN��~!`�oN�����w}��Ů��(�w9��4T�:YaP��y� ���`j�RUV3b��ʲz�,JQ�??n��S����­���D���ovV�F�.�X��a��U�kr�G鄟ͨ:����v*�}����ڔ؇��T��H��ާ�������e��/�U5��z�I�����4T��V�����Y�}[�����
�8Hq��t3_j�eS�p(kTҹ/ۥ���V��E�,�6����<5�?W�C�V��R��xBݳ���?�1���r/5��5m$G�$�C}�z p@����	ģQ͂�Y��e뚂$W�1����9V�4d&�[���1��*(��|�q2��	�?�.��ro��y5d��[^�_)���`��L�τ�Z�%�Qe���5,��Z�>��W#��]��ZJ�ĻF��=d��� 4Q��v��Q�ƍy�����d�h-�y�/.�����lD�d���;��1�l_>|Cg~9��_�$z�F����i"<5ݢx�N �G�8�e�<�d�S��d#�"��[�lnGJ��V���`������2{M�{�[v��-��/���h�8S�#_��P�*���rt>li=��m$���� ���{�c�Ly�H=���y��,D�������`�T&n��ݤ��� ��H�-UU�g���0���ܵ�>����Ӄ��_W��i:����k ����.�T���ƭ7����6j��|X��Y$���<��v�o�'z�Tl��\�vF�Wp�E(�p��/���dX�b��;���[K��^۽���x>ifW��BG����ӚM6��h25��(Ա�{\?�;��\�o���;��4f]�!Ke
Շj�=�˅?��ZK���?�+��)�9�7����ßM�'N���ܵ~���;�t3�0�JTl�n#�n�~W�� j����b���⒜3���Ӄ���@js��&\�D:i҈���DL���K�Ѐ�6��-����e2�w��(�����]A����[0K��7�~ǽ���@�j�(m������M�z,�Sq�#��K�Q���N�ɐx���UVS?
j�k�Ԩea�w�{4A>���5v��Q��TeĀn'��Z����N~�۶�˙
 �S9��M̝����P�KT���Sc�߱Ё��EV|���c(����ؿU\�����6Ã$�u`=	S4�}��j?oA���|��[ܰy�JIq\�ҖI���S���8i���$��`���Qj���ci@��2��y]=ܸ�߅ߗ�M-+����`�0Ǹ�3P7�j|ox�{V��i���Z1�	�Mg�X�<�}�� \!������c9	���s36��K��j� مw��$�5C��/�wq]�kpF��vK4��m��a(�8�G���.LRFuH~~��&��r�<���2���1�Ԕ<̟0��|����\��)�ln�Z�%y���|gۚΞwu�DPibڕG��A��r�7C���S���q���CKgo�.��^	VS�7�O��;�G�q&�c#��9��/1ls�8���
4��Y�?	ԟ[l�P��_�dY2d$AR�6�H�V����lZ
-L��ts35����#?����O
����"��D�t�<��+x�X�16�uչi�k�Vl��j*2�E�Ri�M�O�h�F�qr�A�djу򏉽����b�����)D��9#����d������v�Jzm[S|_O���Bfw�$t j6@�� � CLu
C�H�	�P�K��'���x���"��r(H���?�ȴ�CeNe��&�g���p�m��%V�2^SLR�F�C�����g���>�73��x��9/Ԋ�=I����΍������g��*�������?�#5�����v�Q>����̸�7o����&<al�v�m閿?�qMt7|Y�8��8Q��w��ݓ��ƃX\V���cө�ЉE�X�}^,VS�d����)�Ǳ��eŝ9��6Α��p@�V�m<��Xsw�Y������?e	�7U�,Bt]vJ�X'�Z����t�ҝIJ���0��C��{�>
J�.~���O�|�3�8-��c�9��.����S���'`aOS/
���s���姒ʗH���>�>̞J�p���9�(�`,����5TP���8
�;`���Wo$�*N����Z�ř�ru����4u��̡�[cu�!��O�en�s�_O��k��#>������5��]���3Y���A��N�ݥ�>��nz���p�<��˳��y���a	���k���5�	Ѳ2�j��,�)�-yh����П��N�=>N0k�ߓO�)K������	]"9��IA�}���Paݚ��>B����e""9ի��ibA��L <�!r6�`��Xt�p9�C���0�}��C��`xq�w���BwI�G�@�u���؉D�-��5(���al�U;O���EoFn�f0�*\��(W{��vT�m��:�@3�B�sGyh����EղF�^N���|�~�6�;���(��[�Լy�{O:��*(��6j��\,�D��
"��}
bϲ����0�4���[���´��~Ic�����݌�	F�1iyd�ڸ�-�����Z�a���\��(����g�bϯ����Dn����CU��t�9e`h`VYŶ�x2<���`�O~KɿU*+i�F��(U�^ ��hQ��!W�����Ufިg��p���sUfi�b0����Q���Иy�%d�y��.`�>]�n�-FalS| ��Z�M�%
o�(cH�z��[b�\���\V��۶��{�C�6a�������'�Y,�a��Ӑ1��}-�$G�&�����V ������/T��4b 1h2�G�Ш�VnΊ3��8F�Z��,����b3e.��r{W_et�m�Z��)�O���5��P���*�غ�u�"P#mC\�E��T��[I'/��Z��`�$��4̘�_�
��W�K���o��Ǎ�c���2`{�������j�s��a�z�LL�r�eI�[�'�Q�p�gâ��B]��A�s�!�c˅�l�j�&≳.��6
��,�R��c��"���F�j@��b��4�;��}���OC���o;-�)d0��C�i�\$|+")������L�O���h`X��ej������ኚs�}%KES��(V��j3>F.-^ˀꯎl`��Wq���򯢉'�����٧Z[��ЅI�>�'�^#�x��xGiD��U���}LVf����M@�Z��^:���yO�=��}�W���Z�-�x��4�� 2�7E8seHײ<d Yˌ��d��i ρ�LxO�n@<��8?���:
پ}��4��+r�#X>�2<t����7�����R1� z w5֜�6`��js`�$�������]��w��z���]�U�REj9�p��o���mTu?7Sefj�K�<�1����v�q�U?�c���{�M�3�����҃ꢒ#�zA��W:�$ �3=�'��L��Cꢲ�l:�J��=�����l ܢ��Bl���KiT�bcvt8���ť^{W���͖�^��s��/o���*6uR��F�ێK� �Ɉ�&��5� ��sȿ��C�y���/<�3d�ym�m���I{%A��C�o�Z��/&?˹"%�M9
&���=�o2�9��]Q�D��H�p0��K@�-,�v���t �1V�x~{�b�?/�����Ռ5*7�� ��yx��ob)0�?I,ϙ	�}PN^�������Y�? N��+�=���~axih.��ޛ�N�������ߗ�ཀྵ`�c�F'�O���.@�S+C�L�^2��y��^4y.�濗�|ng��3�s
D��ݛ"+�[�I\)m0T~28~�ơ�%8�0e5�L�t�i���k�>�2�v]<*9�O���B��[ޮ��YYM6��c��X�ӈ���ehVzV%(I�j�S����"
�m�u���EG<[)��Y��/D.9��+	Zվ�z��8��VA���I�pbx�c���&��'��I��pF�~���ؠA-�O���~7�ʔ%G����w�r�f*�@DkAj���o!,� W���E�]\w�'}br�KOR�wx���,y�HͲg��^�H)om���d�9�V�w*v��u=%��%��?jG��Q'J0\nK[w�����,Y�ev��K�t�]�Ue��M��b�0�:b-$*�V��
^ߌ��=�~�s�Ji��`�B���s_��G��t<E�ƪ8��hTgH斎3b�K���)��Dx���ϿE�[�k������S���� ������"�$������Ѱ*�}��c�ޣ�d��g6��ގQ�̃c#۱�:���Q���|����꺺�x�{<����>�RzY���)$^����ڲ���=����?.Ѩ<@>��&KS����,�r�E������ZϽ��8������I�����מxx_��I����묇wt3#�)�^|��SS��UfP/���b�a���)����[��]c��f�$��QU&Y���g�Z�2��?W�����C0�|b����-�F�b��v�.���;B�}��B`����M��qԵ�GB�\z#�A���Z���n��������d���{ށ�ɉ�gEY�X�3~�U'��]�B̷��02���^�!J�e�!���$�؍�t���3�4���oZ�ܶ�p�"�����h  ~��g�L�N������Q�_��&��ҩ?mB ,&Uw�z%���N��z������=��G��Ї���!��/�d�3Z�����(��⻆�pnTjgx�M�g�Ԍ�G 9Kf寯����d�w��]�ď����%��	�~}(R���8CzZfꃇ&�[�y�А��{s�5������R����A�0>�@ඪW|��W�C5�ӊ�u��qg�?R�*�r������K�U�M��ݴ��ۆt�������lq�������>��e"�>x�s(�p�9L�Q5aP�s��Zp:j%55v�@MA�oS#S	+,�������!g��%{�8�Ѥ��a6���g;6}�f�ǜ����w����$Q�%z� �|,F&-��N��[_���x�V��>)\D0\=���qc�X���]k¬���koܦc͋������A�$�A��/�ʍ�A�p�.T����?HZ5��3}�`{�\��S��cD�س��V�Ȑ�Od�i��tm�6�ک�w�����x�ӝ96�7�]ϰ/���LHi����0'i�VF�O�R`l����ī�8�ٸ�[����6����� ��
�f�$,Ѯ�����)ٙ�J��s]->3���N��x�k��
�x�IJZvj�T�N˄ks�PL3��Kr�3}�	�L ��F��ܶg����sÀ�lS�g�	!{R� R�(�Аʛ�m�B;�-�"�\�<����;B��<�̙�y
O��Z%�sq�C��@j��v�h�G���sh`ǧ�Qo�} ��hC��3���.���a�E/��S���m%_��ҒW�E�J��|�r�W���~�-�5{��PnX*��e]4P�����>"���Ɇ�1�١�ⲝ�ӕfa<���O�w��"�%|���;��T���!��P�O�~	Q��m�,����,�%&�+Ŝ�=��5�[/��S�$^Zqr�B�1-�s�)��o���z��HR�<��K
�p�3¥��n`�ȫoY���>��,�K�Æ��f�D���l�c���x�����ip�� ;�����"�M9�#�����k�/��d%>�^N�J����\ hψ��X��)�vVP�*�3Vpk���E�U�e���L�x��d�ȃZm�#mn��[źg�G0�j{��41���� 㬫��ҧ0 �De�J��@�&�r(�I���,�D�v+A���~岉,�⾂]���(?Y_P�ޥ��DU[�Ǿ�?�8���t�>�6LLJ5N��^��s�"6O��1(h��#OJ%����\���-����� B�@����έ_��0=��u�i$�t��o��v7�o���L�Ya��i�uR���Y��ӎr8�twW�a*���-ҭ����V��5>����u�}�V#�h�k�#ؔ�ݬ;��T�ֿ�����3Yz(���;���`\w.ܾcg��ߟE쫖�\F&Ju�Y�x�Xm�+,b�5dGs�����Im.Bt�n�n^(P��?�%Dr�e�#J�ST4}Z��H�Y?G{�b�4�>ǝa�'��m���B`����G�m�սbc�T���|�4�*v(+6G�͉;��1z�v&$B%O��/���[r:��w�d(�"� �s�(���a@�ϝ^�~I�ĩ������貈�bl.y}�s�y�v�𖏫�ק�Av�G���2,��X]��S��+;~�f#q��J)0=c��xt����խ��JQ�灜f����"S�_�nHvGd���<��/�L1蘫0  Ț��&�����ö�7��U7@�!Ar��y��n��Q2���U� �/���
j�b��k|?�0i4��0ea鏥���I��v�~0�� P�U���'�EP�N���??\f���U�m�>������'_J�%� �g��dHQ�Bdf�h�)YY�k�x&L����
�Y�~�L�TBs�h_�>T���k�o�hvH`h9�W�z���̡��i��Z�6�e��Yɛ���0Y�CA���e䥡�f�a1UuK1�EnB|H�$<��ɪIc�g�}(>W�<@o�E�m�z}�|��Uu��-r��{y�L��ܿ�)�7\����%iU��Z��@��4���A���/�Yu�JW�9�W�ˑW��,4������]��u���N��lcZ�L��J���%1\^�mb�q�
�qY"�DT|&�i��GC���2�C��}�^�rZ�e�6;�x�?Y����Č^�-t4 ������ۂ��e�w>s���Ą��2쑽R����`���O��J��7�Q�	he�~�4)/&�s���ܓt/�����Ç�;�l�}:�9YG������m����Pݷ�t�W��͟�l
`_��Л)9P�O�x7�' 6�����u�tJ��35�<�*��V��x[������O<n��3*�:!��>�@ą�X��>R�<��� I�~~�3a'B٤����f�*�-����&7ٝl{
��=��1O��*̴��@Z�c.v*^җ��\�����x0|i�=aX�V�*�W�{�H��Q��K=X��W�ҧ���������� �ci���ت�瘙��6����H( 
7��OW����Z[��?��>�ҷ�l��Z^��v%X���Cji:��0Q��Ă	RK�Y�{� �"T� Z�Q05k>Wp[^b��.N��^�;��,�O�T�]��0M�x_�8��z���i��P��f��޸� H0:Z@ʹ��/��!�1]��@�Gd�G�Y1��j�k�tЦȦh�C��@���W%��Q8�:���<����~u�n�铰��"|�����VnB &�T��@S�F�Qɕ���v�ꫭ�y�*�����Q/�4H_�~0�<J��r3�)�{�}=�~�����Ͳ�c�?�qZ�U?æ4Q�ڏ�蔋x���2i/�?�y�[���1϶N��9M����;���D���~�-�˸�`���CJXJ�S��ǹ�o�iz�i �p+��>��T��<���Ia�}��;J�N�_	8�������Ɋ���������l$�,X�̞�����ˍ*�MM�Q��3� �I��'��ܭZ�qם8�XlFy0G�0�ְ�z�H� �SF��Ѫ��я;����\��5=�ϝh�� ,˴��L�0�����,x1t� `���6�M
����X9ؤ�
Z���vim�Da`M�%��.pt��f�D������vx��~>5e�TF�g���6N�����fu���<s���@ZL�X��G`�f��8��MA�J�y7�̤�Y
G{+
�wS�[:���O��f������������@$l�h��N�I+��UJ�c�9�p� ����`��^�%o���"���_����̮#Op����<\Yt�@s�w�U�Z��Jy����J)U޹��uŲ��P���l;���%��d�
�X�����_q�L�2�����@p�̃�R(i�dB�Y����@�D�ґ��0M�DS�-�=��'��!���T?]�5J7� 4�ìx�k�'��RR$��I����@��O?�&+��
A�
�Uux(�h�б�/v	t�g_˩^�)�Y��s+5�.Z ������T�(DG�M��׭�R�G�U�K<���Cp���%�u��pҤa[i2���w!+zMJ��%q����a�Щ7��GH�F���	E_P����|���F��j�!�����
ѳ}���5��# X�D�d�-���=��2bϓ5麺�9/�%��ӱ2'�y��M��}}�W��˷L����΍~�jg��,L��#<Q�4s�������r ���X��O�$�b�?��~�MdoC�S]?0u(�G����2���C�$U2�u�O�o��I��Ӂ�""N9����C�f_���
��OQ��&싫�)Ӆ��D���4��ʩk&6JQDVn��l�bCp�'X�^��(�o���/ӧ�w��'���,>���	=@�@��q�$n��q�� �_�8�P/�ՠu_��-��7�5�bC��9����R��|���s�F�?8l筵sLx��HP�w�$g�Z�G�E�B�/���r�Y��`��5d�b����7��$�x�)mq�8)�(Hk�x.-7��;�L~�֎���}@��CO�F���x<�����8S��l%NX=�O���H��U��n��a
�+�$ָ�j���r���u�.W?�-�w9CZ�雌\ô��K��
1G�h��Sƾ�k��:����,ˋ��Ȝ�W�gȉ T*���� ���J}|�V	4玧�S%�3�牒�X>ʢ��xW�������P�eV�eA��M�3�'aJ�5tk��F?�ȿ��Xe�l�X�\��������!V���:�,��Y{TN�pNm��{.�)�1�NQ꺓]n"v�����O�C�_��(��e�C7s�ؿ�@�Ye6v�c��$�JZ�~}Zp�g#��:#o&����n�B
L������:>��pX>����@;gv�'e)�h�ּy�e9o�6�L*J�Ɂ�B7A�	v|M��� �m��|���a@��S��rn#b�]�+;�:�9�Ĩ��:��=|݉X1
�
��=����Q4���S$���04��JP٢��7�B���_��Ru%0|��Y^[�fW�6�Ԉu��2;��qsw[m�E}�C]X?
O�nH�7��D�&���������8����~�0���f+�nEhݝ�~ēѧ��-�
��ھAOw���vq���2��׸���/?�� t��LI����Ce}ɜ��n��L[�x�����s���<|��<+��@�n�i���1*'�����������Z9(cU*䁲�t�?�J}��y����Vp-.K���_V�2p)`����8��f=|hr���?ŽފD(|�Y4���$�kZ��y���<���+��5e�CGY(Д�\�� \BՁfD�=t�N�r�v!-���/CC�i�Y�:(l�{z
�#�͍Ԍ��&E���Xn��/r�3�_��m�k�7���F	�S�竽IJ%�����t*�r�L�j���3n(����K�`I�R�:�����M<�����D��G�OI����N��z�U87����Zt%�B�j���4��� ��U�MI݋��5klq;	�8�<zð�6)�xT�ذŚ�����]��(��D�8�ީ{tp�ohT�������߭\�"�6�x�����YdB V�  n �`�[<�wj(�V˰C-���^�*v�Yｽ���$��ے�#-�Z�Z ���%�d���1�Y>ny}��L�B2^8N#�ݲ����#�LF�Ţ���k���jm;׼�nWj�G�N�GȎ5YTav=,D���<AI-�h �lPOR+��$�t�=P��oZN��xdO}g����71Lt��LHK�FR	�}p�ʼ@�x��=;��(U"�5����������Q��.pY��G�yh���"��0v�܂ ������qW��w0��~�*�s�L�/URQM�e�j��,U��3{�i������~5U�8N�� ��Ώ��wު���w/SG��L��̸��A`�@���=8B>��>�,4����+�HHY���3�����h�DK�Ь`4����/I�fwg"�%���c7$G�-�*r�%�J��;n��S�dBe) {,7����~r��DO-cæ���ΡEV���H/OK	���&x�΋Iz��#��WF�j'����#�ԏ=����#DI����40�O���F~L�����ao��=��H�˂<�@I��� -�"���T�mU��3'�:�=�ٍ]Y�Aע�b�g/�794Up��k11��X�����Ȗ�δ�G���`��u������S��jn������h@��@F�S�Á	6΢ܘ�j�m�4�ャ��N��9�@�5�l,�9���~
��9�D�f4�H��5ЫZ.3Y:L���4��h�� L��I��X��t���z#Cj@����%��mO�I2�V/�'x�.?���U$��W7�r�����9֤�Oñ2�^�Z��zlt�N��!m� �VA?���pyq����$*WEd��h�4�y�� ��<��4[�ǯ���E��:4���2�#����B��e���"e��p����( ��a����]N\l�ae���.p/�V�슽���E��!$������ʹ�;�-_�`	�?ڳ�����_*|}z<�b�~RB��<���k+��k�A���)b6�e30i�o�mV6�C�(��B)�*�W�rk*��`B)h���ɁX˫ c\i����MZ��JmU�DsA�:�7�V�A2��I�����_��t��}�y$V�:)�e�Ã3�l�3�Ӆ�r&K��.�)}_͊�����B+g��/{*�y�=���['�L\��Y��5��Țm�w�v֖��Щ���<B)E>���g��Q�M��LZ|z�M�,��Վ���w�m��5���sp`s�3mKP`��t/��`bq�l;yI����v��� i���^����(B�٩�Z6�	��wϵL V��v����׃��T� 9S*S�9�Iv�����N��~4 1qfT�e���_�6�<g�B�ѦVYB9�}�ަ ����9�!�e>{'�~޵j�2$
��w�o��M��!��I���q3�ȍ҂�����:�j���j��Z���U���*���G��z�$4���=Z~��Y��`5e�ٹ"AO��M%�=��6��v��5��WcC�m#������'�Ea:��@�QA`f4����֖bU	q���I�L��e�z'2D�m2�}wXCnmoj�L`���	�y%N��O�W&�T� ��<W$�znϡ���=�.�6�/.�~����Kf�+�c0t�S�"J�E��� 걝7�Ib2+#��-t(@���0=�< u�BV�_���Ҁ8� ����}�"�}�PoS���&J۵�[����f�D3���P�r ��1Wл�z�W��@��ؒ�=�q����u��m���(�(lQ�X%�R�&�Ŷ# l`f�U'���o���F���C���t�-�+馦��~2�?�Q���y�+,H���&��\���'�׹*����A�`�w(�<��;jQg��<-�X�Zl�����B��w����VPyөǎ&tT���}6�M�V�z$1��]��a$�Rr �崳��{*`����V�]**���?�W�q?}�KF|�%�~�����wn�"2k$v��87�Ĝ~}8R�&�4�ӱ���p�����yRe�>z&`/�������u�*�C�[&5�OB��@JH�K4�ܩ���o�\{��ؼ����וX�3�!Q����.p|�p�t�ْ1�xt��`��J4�B&A��
2^G<�����.���G�����&�4>kc�(�<?���S�vd�F'��#������2,��Fo�
]�H�x�PEePG<�g����&���������?L��A��.(H�5͊Y�S�g��P��9=���;y(Q�#�5�i��}5z	�Qe��AI�k�c9tyð8�xy��V�Sѻwp��[>r@��+��;����Ϛ�j�o�@M���_�����>o���'��rP����nt=���m�M;�A�I���_T{O�o��:��+�<��i� �iV���S�|�|��;��<��� �,tY�{σ�(�g��m����%���ŘFړ#��7�/?�pl8h��³��p��ޖl�� hҕ4�j^�<�77:�[��������c����$V@C�l���hX))i
�L(�}��*����}ي�nb��1�P-��ӳ�ڂ��x@���/�"\�]�SE���EZQh1	���� �@s+�3T��a��خ��g1\����pJ�G�!�b(���?4d��I��foKm�̬��I<]������~�E��K7W��k�F�
�Ҋ��;�b�ѓTy.m������;�K�����<��ƶQ�f���	IF6'����T���M������a�w37Y1����h���z#ջH�̛������F�h�\<��0� 1�.A�*�7���v�O��/���H=�B�M���JR���]{x�2�QTj����2^Q*���5H'�ơ48k��>�b�YO��Z`^�]([�h'�,����ʯh�)���<�����gc�0���7�bG�����{e(9y{dJ�z7�c�;7������;���s��M�ͮ�5��� ��4����V����i!Xj�m��fB��W��
_>��7YA�হ'i���-�q����,��P��V�a�V�E����><�V4F�Dރ*s�u�G��F`G5�/ 1�T�a�B���Y*g3��R=��!�~�U�_�N�9�̫]����e_<�bR����h����'DƔ��%g~W� �� �t��Q�9\j���wL�T�Ǣ����2���R�FZW'��*R��R����=*�Eqě]"��!�H�ɦ[mdm�Ǯl���\��<p�L��e�p ۄ4�jp<a�>��.I�r ^l/��\�2�>P61h��jh젇Gn�S}j����ф�5Y�#:���97l���<��% r�+�T� i�%��p&+���<��6�c�8E(L��y�| E*{<�ؗ:�@�Ȉ_;���9d֔t�mWũl��&a}���L�3���1M�m��ie������k�
��T谁�6j�H$_k���)l
�N�r�M�SبA�t�����豂�#�8���Cb����0R���D�#2����Q|ETAHي��� i�Kp�ߺbU�tZ}�D[*.� ����2kc���0~����6e\���h9��m;|F�`��;U���k���~�q�C¡�C��õ�� �m�;_��Ҭ���y�]2������=o]�����2.��dd�;��j�����B���d$y=�����wL�s�H��S`&~Fe=�е�M����ߑD|���?�X_2o4dԒ8ĭ��ˣ}�ۛ��`�TT\0�7������N�_=���~!����C�Z�F�7Y�+�����ݰ(��	������תIU�pCmJP�N��S���u��?ס^�۽�J>�������8S�Ċ��29xr�6���OZ���f
��'h�Dܾ��Ģ@��={G�`�h5+�l�ُ�)��2Xol���~6�"o�}q
��� ����*���x�>���' ���^��a쏾�zQ-����y�F�����ݯlt{�/.��J��.d�mGlq�_}��Ad98��.������Asz��-��t9����^o&&�(�Ѻ��K�MFgT��ߥ�XN֝�	�늍a6R�剫��J{)���9õ�q�T.�?�=CԶ��xωK��|���stk��.O�Ԡg����#�O�zWw���3O�:�5}�1����)���&�_=�3H;|� < r�]�Z}������,p�=����^�X���X�-�,�Lٳ�0���k��M�\��=��iz\s���O��c�N���*fs���������Y�[�7���Ɖ�؝��c���ۅ&o#��C������,V���w�2qU��DiO�fBv�LH{�R������U��v�����Z&bG��"m�����E $��S�X|{�� �4��m���(��
Y����UM�&XY�fӡ��ag�2Z:o�g��\@�2�c �2������CҬ[=�|�-��j���ғ��J,��/Q��C�4N��R�'x��jB0��P
�ނ����x��3R�<����O7A=pO��"�����_|ܞ�u���~L�����o߬�l������U�K<��Rs@lnT.F���ɠNq"jE��W>�Q�Z�1u+J� �Xb��y�x�s��AM`�s}^��̶�覭MP��k�8��f��}��$H����������f+��tt�N��G������:F|�I����m���\�t]&D�f��+�FymD[�v=�nQ���خ���b�-�S���W?w�{��@z�O�B�fs��D��^����r-�������,7����L�?�DM|K�
�Z�_s��g��/���_۝xo���u}w&S���ŋc:���e��箤�9�ĈR�s#~��*;��#^E�*�K�Y���L�l��JFo�.��t�H�X��'N��Ĥ�ũ��GV�6�n���;N'��v갹=+��R����]N���t��źeR�������~�O#�7��|-+���ͱ$�������t\���&(�|�XG~��-25=�ć�	����5{�8��<iW�B�4���u4��N@ٞ�,Ь�P��!#����^y��-�Th�Z~���؊:�X�t���0ηKNB����	��c���e��_-$Ұ�JA�P���ftY����s`��9���X����K�Q(�In.>�Q_*����	4POڜ�Gm���yܵsܵ'���ͱ9��sm�l.�C3�"K�ܳ�|�a�p�l�q�NV�l#�x�'�k�N�U����W��~7�����������궊�Y#����V��͞ݒ��FȚ��L^&�:�I�u��f�����r�t\�k��K7����D���2�j+݇ޗ�<KJE��9Ni��G	��V�FD�Y��:>��ɝ��MT�EA��ʋ(j�W�XU;���q�)�Gn�&(K�ţ�]�2J�b�
�"Pݬ~�l�w�Z�Ҥ_�6"��emyN
c��������{p�Uf\a�-�^L�L���s���&_�dƏ���*Mf�j\��7�8�k[������%�'��d��KS�n^�G��4��46��J����a�7f��(pp�ݥ�H�N�.�e��lue!\k����D���Hd���{��z��X�h�8�R�i�5��N��iև�m���W�UL�[-5t�b���GwX`W��楇}��V��Ok���r�0`c%�j���|5�_��@�X_��c��A�4��n��}G���ކZ�s���nw�ۓ��f羙��j}��j���1�J�ʳ��]�	���*���PF����k۾��ηC�Z�x��}�Iv-�S'�(������߷`���V��P�$m���L�S�v�ǧ�̡D0݇��n~���xR��˲�������ֵt���u��^֛�a�\��N_�)<�m��ʠkMK��0��>l9���$@������,���s�N!�����+${(���M�JJ���ύ$π��3����6�8���s����P�O�%������������ґ�����GIИ����P��k}�A�\�M�e1�n����{!��<�q�&�	7�3.�MT�:�:0KI�]��YARv�ضZBHm�.�.!� M�l��������)�Dx��<�0���VS=a�����<P��}.V�ؽ��������i��ڗ���w���_�� ���$O-ϐO���0`Fv�����dl��֞��1Ǻ&rE�E'5��/߃�$��O��[�
��Y�3l����	}�VL]���DF�O����Ӈ[��0h�L�OI"�p���'�M�ׂ�C=��C�(�X�n/�)��v3J�d���C$\�E�;���;�ݧNd��^.x�N=t}�3�NziJJ�̎��mk��"�eπ��)/��Fh�E�4V�� |����g���z�-\4���I���:�)�(,�ìSS�ؾ{ @�d-���y�T�|������#�u1�	������R��x���nQ=3�㺞ݗ���J��I�����lȖzT�[���j_(��/�W;��E�ʞ�-�گ`T��T�o7��1�c���REGU*��U�6��%H|d8��K8+U���B��w�?�̹�v;1
b�$�30�W�|+�~8��Rs��暣��Ӗ#s�'��:��z=�阐7�Bк����x���aBI�/���a�kv��e�x� ���*=[�X2��ի����J���O'�I�E�b6��*hA9����n�!��5�t�Y:�Hke�NЮ9��n|Ju��"�F���(��1�������0�۽}��&W�ɿ������{��o}����ٛ5I��\6�I�(1��S';��u��"�ź�3Y�-�5�� �+?X:�b��(b����^���}B�2�2�0H�'^/[%2=��b-_�G�0mQ��A��9O�>���D.]]nԼH��U���H�
=��n���V������t<����#¥��E�>_h������I�娍�_4��WI@Z���#��D��?���&?�~x{��Np/�A�x�.���w���ʜ�9��/$��VSP�� ���s(��hg<Y=�ZFԿ�S�|卟R믪�8=+��C^�M��������Q�,��г}����;���>`�����ln_�ji֍��h�@	
Z���LT���ڎ|���Ҳ�DF�_�TY����Y?e1[���#_���S.�<��L�FS�UG�Z��d"W�t�ָ���Z�=���V�e��������~�z��aj���:�G�y�����32,�Cp��Ǵ&�z���XUo Si�»aC�y����.�z,����k�e���5�,��bh�:�i�SK�/ޭ(����uuD_s���Г�?���"+x���-[���5�Ѻ��y�C��Q���[�|q��Cl� I�\�2�����������z�?
���)q�N��܍3�Q����=_7�UrS�|��u��$�%!�h�Ry�k!C��u�K�����x�g����u6>kMݐ��ɹk��Y�b�mo�k�%��/ �/_��/K���{!Z/,��9f���Y=�u���l@��	�����M¡����sbA�s;���O��?K�J��HK+�u8��b�N��$��qޡ��;�ʇ
[i\�;V�N���>�Q>7�T�A��@$��&�\q~ѡ�>`�Y������^�A���d���:�����|�?.�҆u��l�d���=1�V�dB����w=��y��D�s�5:H��_`(c�?6��C;h�D�6mQ%?�3��8��)M��91��q5l[��)���b�5P��;�-�a��[iLdm�z�@H35��@vy�~�^��?���@أa?��d�=�a:Bpdڱ�ii���Ndpua�M;AcJbC�p�Rx� ���~@-?�Ψ���X��o'9g���,���Q9�_��[s����vئ&�b�'p��Ga����W����fx�y3�jP�&Q���F�f��f�Y�2A!�a��|�|ˋ.3���Lz�V��qfT&&�h������{�r�#l��;(������и@�
��x}:�)�tk���p ٗ5�|��z�+���_,��\�ܟ�����9�PUe��j[䱼�Q�T6��孨���LH���a���!�������E����v�6*�fn��gC�ã�%Α���P{�ר�<ڝe�+=��K?в�:�E�Ƚ�{���ds�G��)�E���K��g ����H�X�
E�T�b�S��!����K��RRU����4'�T��d>���mJtg,�Õ�ذ�*��_i]nʉ���N
7��M����0'�u��͓���N,�d��n� K9 ��W�� ����RoX:R͙o�*�?h
��}y�-�b/�Qr2<��=�[��KR�֩7�g[q��qY���GK��D��(�O���.؆ U�2>93��������j��t��]�!o����g����:0(5��U���}��;�{�Iz6�g�J �+�-K���� ��WB�B̏#ߝn%�UI~�:�pR�r"�1La����HZ�s�a�ǳ
h�zv�o)��6Ð��pA��z��\���:��H��+�V^i�a��U��iu5h\M#V��>��#v�\���h��E�����Z qF n����������v��S[���3��ೌ���5��ڮ�w�4�4[
�Ë��.s_�m���iz��t��yg�g�q���ˁ�	���IC;KϮp��}p������W=g=		�t2������k!��#��8Oe�ݼE	R'�A�Y&�{ 6.�-c���?��1|��!�{�����ؽI����OO�1��UK���4��B���V�q����P�zo������*�'�j��/d����tS�� ��?����R��V�{�)���<�|�\Ͽ%/���s��k���+�������S��?5LR��MH,Vڼ����V������k��J��I~~�;���1.n����c?����O�V�_��zi��0w����e����J���v\���Ȉ�#�$�g�L���m��o�5Kr&|�����7$_%Z�)CVu���3�x;�>��K��a7��}YƝ���8��d>�x�y�6ުH�����8��0U���5�����1/�0�P����_��2� L�Y�E�	4���o�pKr�X�/x���B�dJ^Ux��x!򫀈R��G9�����hפ{V�H��r���S��u�z�a~����Ayy�q�9��"ߌ�^����������[�b��(`��AdUH_���i_CyJ�DeE;XW��ѧs���� ��[�8/s�ȷļ�����*�YA`����,t_s_��D��D��&>t�7jfx��I�� ��0@�@��v9���%��a^��/�,O)�K[����z1r�Ϩ�Q�j2C���+-Kw=SR��Rr|�ݵ�#^�����d�F��<�evE���"�{6׀!y`|:���w���y��I�h�c��M�D�@
��䄪Uk{ ��Ϩ�k���V��,�9	�_�a�y�/W6/m�4kW>��M,E�U���$d�,<��A��02Z`����\é'F�����
5�|��#	����:.��
Zh=*���l����P��)k�)�ҽ�f��ѕr�ʱIg�Rh�P����=�`LA�?�"-�{LDP.���]Ø�Ed/q"�����K�em��S�"���8	�ɽbP3����K
��aqO���4��?:����{Wڎ3��0�|IS������b��J� ��=���Ԝo���݄��g �/�0󃋰�!g%�4��Eh��;3�$��Ȥc�'��7u��#�ES�1T+~F��r�fh�O+��%���`�s��x�ŋ����� ����Nq�U��C�Bư�;��q�)� ��9;,�ސ#B��Q#��V��??���-֠dW������PLV��	^rv���q{2�������J�����nH]���$΄����c*w_y_j9@����w�pT�ֵF	��_-<bς��\#'>��O��7�s	��]�`k�
��紡Ǒ����o�<�y[�5#Kيo����xjeSkʂ{��Z�5[��F���vO>�����X�Dn�k�Wj��P�2+��e���`aj��*���*"�u_:�8Z�臦�6�bh��%�lF}tx!�������~�	�	q�A������jl�7y�m9}b��m�'G7m����\��'lO���K6���_��M�]7nc�8'�q8��>�\d�7rO���rK�rb��s�@�y�K)J�L�m�����ɨ6l�� )ax�ԟ)�!9R���Ӱ����Ge���hIn�*��Jd^��E>�v�;��N��m��vUf�X?Z*� �%ϲlQ��Wo�Z!X4�q�Sdf<�J�Ws���lx_Q�%����Ժ֡��c������<�=�����ż�\XH���Η��f�kة��z ���(��r9��#��	�������}���	x���͹����!�|��z�s���A��__Cm��_|�.:ݠ ��W"-K���'OI������X��DKR�� f�Nν��5��qH�}�V8�X�|�R�&�o~nr�1��$r�?�0�.ro�������)�׹"�}vQ�4.Y�ƹn��u����-E?�Pϻ&w�}6:�j�sߕ�PR[Ӊ�������v׃�����	�c`��*����`+B���=��N�.��W����檵�qn�B��U�@�ȿB�s��r-��(��G5�eۖ:\2��sF񆎰#�N�����M�i�,���a=�>^����^�#�␝�P}��1wO�j�	��^n�"J�M���g�P!Y��2J�xmW{e�2�Ǻ&CW$�&�
ͪn9i^L�~ڟ�y̔:e!��z:��ŕΪ?���H�,�C&c���dd��y�����6		��/�Pa�t�!��I���MK6��Mfz��lG�_��r���# ql��y�TJ���I����y�j�.�K�n���a6��9���ppu����(���\�pcˑ]9j��;���1�nYF�������U5�{`	v�-4��V�1ժ�$�#$�]��;��W�8E%��%Jgj�#���$��Z�uMa��X�D�&�4�6��A�.���,k��}z�z��$�~Ue�Kb���{��D
@0�d�?+#^{F�=y1��p����>_1�u�tf��`���
����Vk��|
 p�l�=�I�<��V�'f����T���u��?d�43��A(�XzT��[�R��E��3��[[���D�Y`�A�Į2U
���W��$�F)v��041�inf�¼�>�\���0i۲U뻖�'Җ���~:�-@���_�1�bj��V%ۨ�l�Ճ��*v8��(xY�PF���ǑjBE�4�!8q��̧`w���B
J
s��S���<C���/z,��z>v��+������t��N*�������6@�,~�y���C��o ������so�~�sFYbֻ=��L�7�Y� y�~�:˪��^@ �;��\�[FB<1�N?X �4���9@�w��	4h�H�;�0§vƷ���;E�����j�[����#`֤4��<(���Q_*xP4ê���b�)IH�������,@>:cc��_� �/xd����kUp�����e1�?B{>I(.���3htt��az�(��H��NY��¶Y-ҧ`��	S��Pc����w�v�Ȳ�!�릞F�7-J���Y܊�4�*��u�?�T�W|�g�D�u��=ۼ��>7b�I`��%�
���vu��_�婔I��L���q���N)��o�FK<�vK���FK��-{O{_�Ey����_'t��ӏ��C�˂�L��M��mfUF~�!��v��k(x�p�y0��xU���*TT�d��՗-�|��hV>8�������xr� ���&::��H��qp�Ӈt� qF}��6}'Iy�	�e\A����5퓤-`N2�:���ӷ*��"���H�Vhf�~�l랁�Ǒ��z�1~O|���VE�Vo&t]qA�������:�+\�!ڃ8�Px�<�1|HāP峸_���qh�+�9�`8��	�׀o��*  ��Q �Wj�8��'���ܐF��[�|��w���,}���<Ґ*�K�
���&g[��N����^�{���@��g�X��՚�2o(��������f��,4n�?F���ȱ_�K]5"�{��ݥ'�0�m��#쭃�Z��q��)���;��i���������{m8�y�w�ߏ�3s��}ｮ�>���ܥ�ԁ�S�k�6yW���.n% ���Ħr����n�SX�ð�?���A�~����Zsv��ߵ�خ��Q���еK#����X)�Bv̦��S����#N�Cv�)U���|>��������{i���B+�~�x�A�����h�}�=�L�r�9�Ŭ{A�8��b�|�;���;��{��j�v�ob>yx[9��N�`l{�0�����,�	�1����I�qu�P�)�~�XJ�"�g=��)V+�ih'�h��-��q�K�q���L{�C�[!��"�?u��
�O�cU�W��An�L1����w����M�W�G��	R"v<̂ v�ū`�I�!Cf�q�c�ZnE�i�	�}fg�Q���&���>���f4�Pwۑ����g��������L�Ǹ��W˛dK�$-ר�M�{�u7��7��UY�\ҿ1yW�]�ʹp�r�H��'�p�p�=�ܦ�܅���]k󾢬��C�����$�����ޥ�ݏށ#pQ�c,kQ�a3@F�v�5�o0Ͼ�8c}�X?*b
.҆��3��,�dM������'oFr���s]s�ovB��;����C`����T����c��J�~���{��B�oF�\�����H�)�z�<_�L�h�J]��[�|o�Q`�漮�A����e%+�Ѯ�~�=�B��. ( ��Y��,S��j�Wq�d=RR�^N�<!���g��ݍ��%��յ�t*8(���w�h��_J]�J]��9(3��c�;�����u�'A)�z�^�&c��o�71��t����hC��u]�:P0T���|�#oo��J
�MG��_Ӧ�'c��b�h�ˎ�Lhz{Y�d�ʇD����A[�Oܙ�e �j�y�o�^1�+���?oƾ���}5]/�!��-y���$�#+��	ՎIa�y�aC�"��&��E8s���p�\���+�<`-��$����V��)|��?�v���%V[o��|�y_��I*Sk�I�S��@��Z:�j\�uy"Xߢ�$V�+6�������?�9��Bk60��)�+S{������r@ٯ��M��/U��Kɑ@��q�_�	5���7����(7XL椁�����P}��z5�����ҭ��&�^��p��q���G&��$*L٣��G_��~($��q�����?�=��Ȳ����K����Á��cf:s��&-l^�d�x9Wcd�sV0�0��9�jU1���3�C�;���������
�g_�-���.[N���M�/Tq���J�8�E�3	��	�.m!'����i_�v�GA�d6��_�5'UW��
��x�"+r�r�v��۶'3�,�B������dH�V^m��&�M�������y%�6]�9�5������r؍��Tnm\�E��� �w�����)K�$�H/�0�Т՛��7�F�(��\����������uk�5��bj����Lj����P3D��+��뽓Y��?�N�X�r�p�E��y���c/�Gh�~�"�j1����%����<E�.b �0�.Oq%
M�ݶT����e��q&��P���6�v�Z�ok����uJ�2]�Zk(@�,~�nNk�Pn#���,r*�K��$��/�5L���ŗ��Mߠ��k��5�B�-�D�Bx5�����[�d����R�f�C��C��j</����.\�_�/�F�#;�I��mcp�g�� ��PIr�
����Ö�����n��J�G�9��m"8pz�l���t$�Z�KP�3q�_1q[_�wߝg��T�uj���D�W��'in5Ӷ��#Z]9t��X?7O+8k�=>0����ޢy���q��M3��R�(�����Fڟ�p��E�u�G
f�|'C��o��њ����I�O�����,d��#��H�\2_�A5g�n�\�EB0X/]�`p45k�:��*���
�:y�[���d�4���/��J'�ejʥ���@�.��,���%jk4���,�5gn&#�0��mO��5i7bbu���ޒN+$�`�UwG�+_l��p���l�e
�i�0�L�^�l�b���}���# >Mm�!����7�k� ����jG�I�:�B��!�+'k�0�]� ]ڳ~p4+�,`�,ݝ�5*<�y
+����U9S��=�hɷ���m����%��!Lv�h�9��mL��0tv�с�r��
5�w�Z�ݖl���^&C�Za�E��e�9:��2[-�oL��Uc=�MPQ�9N%�k3��"i����#a�{텞��3W(I�֨s�;�̘%
�I��_̥M��d���s�rרY��wJR�.�j�Q ֨�����^��/9X��'��U��X+3�y\�^�cw8����kλ1*�D��b4��g�����ǿ�q��R5�텂�㉬@�ω���`�	W��4p8y���Zm���U���lۇv8��
��R�ҞEk�ӻ����n�7z#<�W��Y����ܷ�TT.;#���6�qڵ�g��?�����G�G�T�6�r1�O�r�ۨ�4b1[�;�h����c���-���ښ�?�Z�
��E�tS/lh�15����� W.�a_s�$�b��f�+��C�h+�n���]%|7L~�<�����Qk�������\Z���5&I;-�&[�'"8�J�@D�����t|�.�����&�I�3�/l�V��a����3���W.>y-��Q��x���v�}Q'��x]�g���Ik���C}������;9����靶���m�G����픫!�
i�ۺ�՟�)���33{��i!n?Խ@'����2��@vd����{ڴ�1P@*���Fc_=��i�y�>r8vC�/}|T��^��0Q�`hl8�����;YfT�W���;8�/5bv�,��e!F��@ݛ|�R^����~��讍#ec�w���םg�>�����G-/?Y �4����@An��BVe&Yg�-�,�ܥp��s?���$��[��.�O8,^����W~���%ٟ[,�ȱ�HE.\St]��Qբ����Ft�o5��u���+#�C�������*�r�j���,�YHy
o�q\Ox�K�|��PoF�R�Þ���O���`���]�٩K���,��FK�0�Y86��-V`�]e���-fe��~��5��Sʨ0�o�Oj^[g�?�ɉ6�������.ZTiٛY�;�H�GY�F/~���I��'P���c]��k@X��z6#�H�F�򄂏|{f��~��%p�^Y����߂o�ޗ8���&Qڽo��ީ.�(v��J� `� ��^^�涢_��@5u�Ux@b���C8L8��_&�P��:��T%bj%�hw�%�x�N�h���<2��;�����y��Z�B[��:/�@�Б�.,V�arp/���XXT���Q��y��,�.ܥG@�i��\$d\���- �_��|�!�:]p��t��M6-;4w�+$��T�;����M�v8O$\d��������[B{׀!��8ʠ$�[�� �G�Q��4��x0��������l��h��q�q�*/����l���K��fc9܃P���
���U����w�m@!�BG��Z� �Gjh&�0<��x�+D�����d-+��r?&Znz�ݰpד^���`�o�M�Bw5��	=U�h��C�y��޺�ug��)�e_"��0�w:6�f�v=}v;0��1�1r�;,1���-�Vjj�_�O����}��-Α���/���1�=��߹�7 xpD/�?2Mb$�mB�� �[I�}q��LhC��wo�ͧ��^ޤ۶m���(�z��C{����
 �Piý�ta�ոX��G��;���8vv1��8

:���Jq�Z�Ѽ=z/i6��fj�6�2֦k��[��:�?4����x��v�����(1'�h�f�*�e��iZ��M�ct������U��A�+R��=g�6��7Os��b�tj?���)��$8-q�9����!�@�����'�0�R�F�w��}ۙ�%d4Dz�����\}-5'�)�}����~����f�c��j�-+��-�dk'��I@K݉�Oo����4*6�ޛL�Oɘ(�{N��V<uՈ���P�=֧�)��h�_֕��Dľ-��G�������xK�_P�/9r]kX�fl=vOԳ;c.���r5b���N� J�Ku3�⒰�\�fZ���U0Z3@��bj���_��D���;�1�.����A׼�������Gm��l8Y�,��P����7��=��^����&��h���pDƬOJȰ���g��yd�(N��(�^}����Ml�"!�<��`�����(�ؓE�NvJv�+��b_�M���#߬�*�u��}�QA�p��*X��n"U�������F�l�SZ��p�r[��T\�j=��ܮj�7U�,%�M���=����2'�o����5�����p,7�o�-zs���D��H�w�w�x�wE��jY����g�Qn-��D���NM�����v�t����]q����-
�+�p�̵��v����~ (����ő�ݨ�_b�	#��~���M5���R�n[��)
+E������������닖[�%Ih�,_��C;bI�'�%|c���a��X��[������~�5|EA���۶�]8:r��狫^	�d���t��մ�v̺��Q���m���;�R�hR�W�[��I�nJQ��H.��[^a.��/��DT|n��7�{��s*��ll�GJ�uX]��.��	��"����˔��Q�.d6HO���q�j�6� mq��]����B���2���P#x���g�6��p�T>H�����*̳��������(g\��-Σ!8@cǈ�� n�Ï��~��A�,���1b��q��:�I�,?(X/�Q�`���j9������<�>)\{cY7
�'�6O���"b y�C��2l�j������~�F�]eu�ӣbƶ�����fõ�OB���(l,l�k����%Gq|�-�IA�;��Lr��v=Wj5s����ڵ��c�"��آl�ԙ�v�[?�[��H�}��o��`^��,)񷽊��;�{�u֮(p���,���yT�[��Q���Qi���56�~B/6���#���	��A4��Y���ʆ�( ��iY*��7�ѫs��O(4*�����5����
����tݪ�a�������|��4^p?9���{ɢ{�FUvEC�"Q�RӀ�d�SaMf�yt�����I�|�̾��!�W -��TPi G�k5\l'\D�ͮ���]���ã�w���{I:�9s�G�[��s�u��9���*w�ת쁼�_���{�x��pO�Y�͡.D[ɬq���AS�Dt�I�.����ŵ-���8+���e�1Tl�=��Z�������:d@�'�ԙ�vC�iOhws�p{�Y�%�>�^�!TC�[��P:�3
�����+�iȃ��cF��R��.f�4�$#�<ԕ5D�a��w��|%L��y���GF���0��FZ�ѡ�ei��t�ms^v�Rn�|6C��g��<�p�Z��L��Q6Un4�\��������QA�9ӗJЀ�f�6P���:��Y���'�<փU�&bP��Fgo��x�#@K}�}M��H�q����V"����C�ڑ�������HI)1���թ&�nV8�������4 �JՐ�u���C&�n5�ŌbZ���!KG1��`���#�V}5�8����A"zM-��p���R��o��et?��j$̙Wl�Uz>8�?���2�.O}��[:z���>YI�~Wl�<���yAP�mnq��J׍�'���􏹕�k�d���d$��%�8C��h}��J#C�ы�<�0=��V�hQ�A�rC�ȯBp�偲�&��d�5�����%&���d��:�S�Z!�v۳2������Bj8*`]�9��WA|��t�	��m��c��ʥ�2�t�V8���Vl@����]���м�A(-l��YB}s�1Se@��[a#���xٯ>���j{M�n���%�gH��P,վA 4�&�.��+6'�A-􎤡�iť&�|j��j���_�Ҹ���}M���!V�V��Q�F��~I�򖕯N!h@Q9��m��B�%��	�`^wB\����v �m�C�ϒ��[��l̳���R��Ů��eq�e�C��+�WE|� yf@��#�1	o�dj����MM&s�Kl=�dM��;�����/?3$z�KC38SP/��ⲋ�����G�)ȳ�|X�6d��h�f\ �����`a�e���˘�{��������˕�5VlOBA�!i�k[��+"ޚ��%�C����}�4~�'��7�7�P�]^v�0hn��D�Ql�\ޢM����xV�����8x�"��(Ph�~q��XK��ҹt�j��0�a/�zb�����h.rԪ�A�j}�Bv���L�B�5������������6�> �M�������]��� ߬?���mcT�}�#�)��1���R W��	�~}��������\�^Q�%�%��м$ʿoHx}���W�J�%��+[���kۦ��tG'�݁�d�4�(�6���q|��LT��l.� �4#-���v���\Vc�_��漵���;J�ftɀ$az����Q.r�F�#�.,�/�h�p��?I͙V
�o�D������;�?��ֱY���G��\�.g
K9�U���ȉ�R�*H0#��\��ݞ�~W���q���v�JH۾j��o�E���}a�4���J]
����� .��|C�.^� ��2q��l��>Z������m�+b�B"���{�<�?�=�w?�G�1I�	��������y�(�&{��w�}������]�!�2���j7*�ڦ<���'���H;zA4拼z[][�A���Q��ݛ��22Hh��7��|?����,>�C�1��4gkJ'�\�=2�3�gBD\T������R��=&�m;⟻l�	�\�:��g�Gښ;�M�b��lI�bȾ28st�l\yl�I��N�R�Qض��k��<9���{n`��/-.���/�0�lq���t��&�A�͚ےLը��Qd#����yc �w���P�P�n9F��YLv�P�����ԽM�q���C��69������$ɩ�0���1�|Y��WK4�p\�[��L���T��LN�,�����{�?�ʕ�ъ�ԯ��J��6��I�^W�}$\�H9~"N����;�J�SG	�;p~��HOH�Ƨ����;Su�u���:����+$	�AD{���k���m{�������xT�k���4��d�j"�t$�˂���}��v�L]�u�Oc����F�'�.��	�;i*e+�)���a�!���
�?m^�u�v`l����U��TįD��7��M�H9Z��/�DR�G'�{��0�Nԯ$�臒�9<Voj��e0>�v>8}��	�5M2�A�ӏ�C��m��ӫl�ha�d嵰U�B�7����:�?��Ka�(����~2������6�V:n{HV�3�E�>V�ƀ�����?�9�_uIFf��5-3|r��������N�0M?���m7�\}y�˺i��HK�I9��y0��8�hc*k	2з����U�\�s�Y��q�&��y�<~�Y�J'���O��!���+G���n@?����
M��6��s'����L�QLa(N	���Ŗ}�q����C�R'"�l����ȯ����6���|_ܓ�\/�t�yS���iD�������(�on��I<5��Tѕ�\F��iN������K/�b<�R��l����8�O�9)"�bk3X  �;�ZQ	���q���Ћ/~�)Gk��{���3��Y���	;�m����6�?m ,%"�su���5�F�����݌ml^Ƀ���M�kng!�8��տ���˿� �ݔ༭�Q�j�:��&���<Xx{�)Z�9\C6��G��'�q����7��]���?i�� ؐ��Xo�y�z�����+pj�G���U��Rp|���'�$?z� {�Gr�Ә����8hǟ ��h��?���M0��kW��o�����z��b��rޤv�BXn>HB�j#��x=a�OF�@Ny^]9j�4��Q�Ɋv�>�;���0�2w%E�D�N��/W�|A���1RÒ;��镲��Y��
k���5���X	�y�q`�#���ɞSk��n�~D��NJ����/}�q(!�g�
o5/�l�Ϙl��/�����ݺ���e=r�r����{�.�Z���u��JlUX�g@K
�s��5��^��{4 Vǳh�ꃢ���+�_E+���0C?<v�3����
�Z��,�@�N�?tzZM���b��jB|?�OjM|�Y��)�r�7Û�0�)�C5ܤio*�889�%��Ց h9�?cf��Xx�Ze��[����g�5�6Q��������T�	7F��B�~�㡳1$~z��b�S��Թ��gz���I����ݎ�j�3���߇�} �F�.[�4��n�1k�ͅ�|O0�	Rt�6�X�M�-�f�~��g�^i��ƚ���O}^i����*�b�Tu�'#�c�
p�]z(~Cc��P,1֤�7��u�?F��Y>�1���&���)��l6a��6 s�����,"6���XxLB����ޤ0Ք�z�+���ɯ|��c��=ۥߎZ���>O/�A������� ���_i�n������S.� �-�E�Wߚx���#��$n����/�[�e.d���,P��.L�T����j�m�g٬ttgOhԉ��<Y���D������LL];�_:3)j�_S��ͷ��!�8�Tw}kJ��s��d�$3"������媛<l�ZD�zp�W�qN��t�W�s,~��};KC�"�M�Q��A���i7)z��	@5�mz֗R�Y��<��'$�Lg��/�[4�))�����=1\��r�4b��H��πft�2HE9:�	�, �
��f& #MyI�%�G(�25��h�|�|Hʜ����;qڷ���E\�̭/����$�������j�7p#d�1���I!�[���_�m�v��W��gp�fg?�=~^�0mv!3�1z�&�R���'g�.B�_�L�9~y�i����N¿kH���P����rG����յa�i5�F^vC�;5K�d��s]6;��7l���%Q)\�����ғЧZ�\��w�xH�"ЏJ��(�UjҪ����D�������*q;>T�#کD��w15P���:��C����/��~;�4G<��A��g� ~�n��+V�{'�M�8�5�u4�sQaỜ2�j���2�����Z����M�.u�������}߹����v��%<Aʒ�������պ�B$������G�{m1fJ���<�c�z�Z����|?	�ј�l��Wbe%h��`o�=C��	$M;���F��q�!��B����79�	�2ʍe�� "����r:O_�g
(�J��hͯ�4񥙘���l��n�}�!Ͳ�����0�/��Y�9^�P�(9N6���+RNm��)N��?��j����QF�����"��7K _B��kòt��Ϳ@ MT{�_sh�6���|��I�qp�O�mi�4O�PhȰ.�ڶ��G���x'��rY����È�In�
�}� �w����3�;p[P��~����|�0W����",l���T�D  %���C��.,���i�S'�/#?��b	�]�G�RyI@Y���åB�q���Az	\����1�f;\=����X0x�jrl8�r�b�pi&o��	�l�v��Z�_"a ��}'K�����8��9W��D`G���E�W�R=n�5
��0;�{��pv�-p�� ����~���t��FFl	f�n�rP��@���>Br�J�<�p�ټf�c�.�H8L�+E��:M}��Pl��f����0�m�ؕB6f	@�r�s/ �j�Up�f��n��vh�;<y �$�m��^����|�ur@ܧ&0�fe����wT�E�"�E����Z��4P��	׌%%Vet>"��XS�ĺ��u:�޹��h+���c����W}�^쾥U���ō*Wz�KW(�:\j�/�(x=����r���פ>#���^�*D$3n�wϖ۾������Љ����ǟ8H_$��k�-M���~�{9�)��!��nno�k+�,�{�W>��ge�]ʵ�X���m�I����{���H�46�z���2:A�q�S��g�jE����GkCu)��K���4�J�}�Å�6fb�(7.�E*�IQG�:�`��O�}�s	���=�g'�с.AC5{N�><X��F5�`6��UHOH+i7!��,�tK���Z�a��SU��0�8]sIn��S��0����u6��"�
��@��j|[�����	��V\�~�C��5!Њ��M�penZ�Qm[|����g�K�^�q_^7�K,�"�3Sn�a�_��e/��']%,CH�F#=[!ϰv��<�k���hYYX
��a(�[���z�F��ATnR��|,LJ�>z��Ց@��m~��Te��T�K#�lm�:޲�Q�Տ[��?�VUf�F����h�Lv,،L%�E�p沑T�PھlKJ�􏽺α��d�����7~)�|Q�s�3
=m݃-rƧB%�!���W��js���u"|5`�ٛ�*R;aH�mf�5�g[[h+�Wk�q�[�Ӄ����?�2����얦b����]�a�3��*!{
�e�fxZ���-��O��bi)�A�|�7�b&8/ȳ�0����9O6(#���=�d��z��*��{�Zz��W8�+���)����?ߊ� ���^Z"��l�7���{˥j �W�?���"��,�0�JK��:�����MI��=�$�R�\�`����֖� #y�.�"qڮ0�E��+�>u"jG�ׄ�����8,�K�wAq�W���}��(�35��`��v,/>f����}J���U��	c�bF9:E�@�eC��o�*�B�]�H��ԑ��ɹ�@#c��	��jR����i��䘭��O+��MW���MUwT�~X����m���/�6�wk�/���I���@����a����*Aƺ��;��l�� B�� �c[[Žs}Yz��Ҿס��l(��R�T���Luj�+�!m�ͫX��7G;�6x���(pu��u����`Vw� ٪|g����ܿ,��I�����qy%��c�#���6\v�s�lX���46��%�o�B��%��_���E#-��~���RŅ,��K��:�@L3`��dƉy`��q�䴁,�y��+qnF�vvs;��֩�f�ힽ�t�j�n�3���"氰�n*Qj��1�)�Ѽ$9��]D(ӆ�d]au��̓����E�Z��o�Cd����C�mHxmUT���ya�k���Ʌ�A�\^@�u�U��71wnF)�+���!�`KRuCe�Du5`0|��!�[�����K :x�P�Pś��ޠ�[UU��1�Q��+Ղ\4Z��A���+)�RY��E�{2 ��#r����!��"m����~���$!:y�B�$7���d+��v�P��=?���&��F���	1���[��+�ڲ��eb�_�H�@�^ �[wf���Տ (Ud?��ũMkJAa����D��\"�6^� ��' �]�1�ؼ��oOޤ��GU�+tS>*:DĻީ�^�!�n�-o�;9"�
|����J���Wg4ԥ*b��UP��#�"�j�{�*�{jn�6�4c��"ԫ��r�����Xz㈄fw�Z��Fv��0*Èf��j�,/��Cc<�|��t���;U�$S�2�� �a���f���(��k_A�~�\�a����!J83 g�7��`�Oj�;8��f�f	9�g4�-0�nXӓ?�;�5���ܵ�=������c��L���[��K�M eW%�����> �o��s>8���Mp1K���Q+,�����/=e`Q��G������G��U�ZOv���^2s��qU�Cx�>hψ:6DabT��4"�����M�D�T�\S�ׄ�{�_w�u��f~�~��0�/�U�=)�Ɵ`���wxI8DȦ��B=�������@�����E��h_�$W�B��=>�s�zYs��$?UJ�b�M��5� �[�f�O޶WF���+Eh⅀,���e��3@��4�v5��v���pkmi�^fXZ�V�!�,D�������W���a�w2������V)��b�>�C�>=;HQ��ݓ���GH���S�5,�1������>	�����w�T�tP�
��a4m��|ݾ�up*6�
��=]���{�JQ��dK� ������I����h"1"P�+��ƛϗf8ƾ-� 呁Q m�/#�X�7yo�� �k��V�J\8��I$�8�o��x_%$��Ou�������j�c8�&s}@�گ��Gr�
\��1{�S�ґ�-aF��kK.F%���BC�n��vb����u�w~c�hmw �T��4�g:��7ȳѯ(�v&�^� o*�jsT�@���m��{�m��H�O�)5��?b)��Z`-����y����ں=2�v�E����Y|�@��4�W�r�	/Ԍ��>$�Z�'#�R��!��yDq����=/1�F��F��9��=`�܌�N@����'U�`�a�NL��Q�Q���Ⱦ&X��E��C�Z1\�����;�W9�t~�\��W�����1������t��7���G~<��
�+,�}�/����B5"V�܆�'�S����n���?���b�2n�K���	AI��ӊ�Q��=2�=��g�'.�7m
���x!Xnsm|R���9��=��ՙ�կa�����J�uW~n�Pm/ ^��J2�����[_ƃ���'�R޴�#�XJd�kr1��$�5i�͟���1�q8��%��>B�NQ�������O��"��g�x��y��!4@[�e�!VmpQ ��	����v��$�����)1\�he/0�������[�Դ_R���z��E�:��ݛƗ�����ib�PLƦ�`�\�i��q8�=f*M2�,�H�G�k�+��)O��
Լ�o���%N÷�q���!Ny�۵���xx�~�
�(/��>�����zR��`�V���J���)V����E��)L�	'c��`:�l�8���dE���9LbDo�S�2	���y����~yd���X��i��w�.ϱ;��=D!}l���<�Xх��w݌M�����gm�lI)�$�||�&�x���L̪�����!FBΩ^��z�`\e��LJG�J�pAˏ��j�f���?
d~ý��D
nf�,�T �_^�3�!B�uҺo�c�X���PÅ�hc \b��$�����ϒ.��S���.�oU����D�Pr"��n��^��'�y���`4m�ιzI����l���D�s*%��x���=M%Ǳz)�{7��4���2���ᬖH�>�5L.�7��s֍�:�fS�	:<�3�`o�����Y�Zk��ՅD�����ɚ[P�RhI>���\�?�h��cGI������~�t=Йh]�� ���i�W���Z3��.����*���Ώ��^���4���z��\8�q�q?���9庀�)�y0�z6�[ۄW���>J,�������Sl�2OF��I�3��w����v�T��O_ц�G��uA��bE�
�*(�n�K�7 �Q�&��\}���mޅ:i(GKUN��6��.[C�|���`JYD�L7cK��$��yb������6��=ndo�PX;#���V?x!�� ��]^{"Xr��B|�������K{�
�?���V��IrЉ<?��������~���'.�-�%/��*X켷�k�Ĭ��";_�{���{;}C��.^�[Y����4����m]
?�nI	��*L�����	(ٷ�xOσO��ML�H��`�=�(�F�{��K�S�q�y��Q�V�a�&���oҨπEq�(���h�"��[K&�
�}�*�_`�f��(�o�w%dɒ�*؊ $���g��JDʩ;?�TD"�9qq���Ɍ��g��_π ���M>8x����X�փ���?L�Z���7Q&XR�8H��h�\���9��a7��",�4��rq���������t.w����ݓ���"!���09j%>2Z��i��B��f��V�>HЙ����|t���<�}���CZ�|]>�4�wga.XB��5��冲?ʘ�\~�S.[��GD�p
h��"��?9�&�E>0\����C��,��
}���b�:��Pt��=���}�Z��/q��v(��G�ǲ�Q?���B�7P�L��Y%��}O��7����� �qvetA��^
T/����1�0M}���n�Z�:]&pu��?$��9�ﶲ�m�Ah�\�W�Q���&���h��Rݴ��\�Rn�G�&�d�q��7�	�þc��&x�7W݁����\�.��L�55����;x���J�@��1	����s�;(� �e��-���ڨ����)�C��gz8=����|��e����aÅ���M\�C�sҒ��:?��8VI��< ��}�I��,HH�F���x�kW�9dB��ަB�	���>:~�Ok=�)	
����\��^YG~�ǋ�'yʊ>U�d�������р�3l�/K:�S�کŹ�X��R�o@�XO��9'�o��]|�G:l|�5�"�R��  �q�ATTō�G2ѝ��-cC��D5��1�/�gz�Z@܋?�@>� ��w8��F�)�������N�*�L+&�4�*���/�g���#f���˸4h�m,���9ѯ������]�73�ett��Ӌ��?��osfA��p�{�':��J3ْܛR�a����]���,�Ze��������<��W�H40�g>��b��'K����_�-�;�!򕖦��/m�\Qb����5��_	͟M$��%\X���]�H�J��VU(�M�x�f�	c��+W>��o<�?��U��f�ҕD�ѳ9V���9�Q�p�l��`l��M�,(�Єɬ(ޣ�{#�<ó�������sfF%ڡ��i������Vcf~���?�3����$&ϴ`@0H�$�Y�s���J��1˒�YR���c꒖�c��{w9�����*i���tj#��d�{��x�(9Fh��u�����7O���q0`�w�$����c�����7�*P�j!�']8��#�p[�:R9վ±v[�?mG��#j�OL{�����<t�"��2}T���#�*.N��bbe�����(�UΟ"/3�����?�~����z8N���%��{��
�&R��f�����J�\�+����X&)3�
m�ނ����cXDT��+�Y*83;���0e�e0���I��T�	/gR=^Ȧ٧\��ӧ��Ŝ	t�n��FL�L�G�q��#Y�ӃhI��8��iΪ^=�GZ���4�4�8+����ZD���*�S�r�!h�1B���\ʇ��s�~�F�rz F�<F�P�o�� <������^Xo�~T���[Il��A��2<���8`צp\W�&UWB=��V�}�]<;�Ŀ9j�M��آ���d*��c�m�w�i����z6P\N=�$� x�w�yx�uj 9�Ѵ9Z�!�H��;���76a��=�:�>�!}�Y|��6�]�@Q����_;]����٨���R@�9 ��.% Y�z���4��g��0��0���U�z&�",-�b���#ˈ}k"D�����B"	�����?iU��7�mO�I�&�G���*���$u�FF(������2C����+`ȇjhK���_�>��b(pB�+�ܧqY�i,����r2��@c%�T���>��i�j6�&��p��=�9�:~l�/%���o ��s���M�C�PZ.�{<�c��qI^h�I���q�>,3��īN�~x�A���W�`���%�Lŀ�8W���7ly��x ;���3��%��
[�s�����̊���7F�E��2/�דmJfF��`����R��ڐ��M%����+�Z�����E5Q���p�,P
$^o���1���[�m�h�Tc�F�^p̂����=d9�-��^�ܬ2�~�,$��=I,POH؟��%�3����
؆ʰ0 �:����\�ܩ��L�/HI(��[u��K�к� -�̗|I�^����P��l�BM�=/c�� ,���S��R%e��&6plY6x��yq���ixD�A�?�y���O�y��Y�O	��y8�̱�5���Grq�H�$�9y�NS�0
V��s>oc2�N����<�
�,��߲ᓚ��C�1��r�3b_nsk��f�P$i����M�s�b-����iW}����{�7*��1J�J����x���T��g`��v�ӊ�+��e���[M�J"z�WU
�R^O���CF�y.�v���k�oSJ.��p��a��3֧�L)y�tz�+��x���-�X�]ދI
�Q�,���5~�o��hs�Lx�%�_����#�Rn$)��-��b���//�A	8��5��_o�Ts�DF�`v{��(�%&����jΗ�p�.?��d�ݛ�J6��7/�� �sO����3�]\�����Pʮ��֋����]:_mX�F�fR�ҏ- ��$�Ѡ�5<{�k�=�r��}�E\��iT��e����si:Q2��
Z�4�Q��#���m� ׯ����j���|�	t����Zh���|����.6�*F�wl^'�,@�<=}�t��O{MN�M׵R�Lt���I'��2gq�K���o�T�Jz��_�}��7a^�P�-%��*C��,|l��x�0
F%6Jzt\ӿ8YB����u/x���>!��Ni�g�lj'x
�HV����iV������4�֒�j,���El�Z'b4"����<�� ,N7B�L��}��� #Eۅ�zA+��΋�,k.����&,�Nt;I�s��g�4���9Ԩ_ǝ/
���-A\��G}rٕ~��d���2o�����:�X����y�H��V1�`�6���D����yq	��E�:NH�1ǈa��M��Ϙ.Qq�G:��S���9 ����X�[���t5?}�����PmˉO��6k^o��_7�9Es��0G���>+�T���	@6����༑�$��a*��_��|�C�{��P�-Y���`������c�G\�foJp�����6#RR��[:��_շ�?��X�H) JJ �%1�tw׈�H7()�tΠH#�3� C�o｟�Ϗ�9��qf���z��������r�t`Z��$!���d�y�_�&�������3�=Pb*0�hq�5����2�u�v�z>7?KuM7������Y��7$���\�F�?��w��B��׽f��d�I�FL�'�(����o���yf݃� �I3-8��ټ��������p�7_V"e���
-y���-/��W_!>� I������ŭE���n����Ʀ�Ɨ��^vn��w~�$�PI'�a�1E���V����
�)�W���I�L��}%Kd�߬�2'K�ஷ����{�L �b)����%�(�I@���OnO6�t&},���}�*ŀ)0�&je�Pt�V���}SI����N�W����aS��G�ƫ/�&6i0�,8��O���GR���I
�O���6�f��2��x��b�I:枨�S f��`G�U�N�Qt�:O�6��3wh'(v��
-(�J������ڦ��!����7�g�u�Gn�{���91�]����s/BzuJf�u0��8�M�J�X���4�51�h.���Y]�����x���鮉�YȐ@ib����t�ף����u��"u��Ǥ�t�u��u]�,"Y��\I^�����M�R�7���M`RӰ�;�D��Ǝ#�0#���|e���e||�Xq ,ff~��<#Sس�J;�b�%���puq�I��*��L�+�R�&���c�����6/_r\����f���.���Nd�� �G�)��]�����EG�&���s`; ��T�̂���.���J��!Н��[��޼|��7�`InU��|J˙��x��٤f<�:E�ѭ�j��Y��M�mr�Q�р���Ԉ$����B���?4}��Ğƕ��;;�(Vcg6��r��Ӿ?�.�^�,�>��M6,i�� ��e�Vt��;��yf[M���?R{G�%3�<I#)E+['���h�ֳ�RG?`!�P����vط��A�t�������mƶ"LBL�dI����!�@�\2���"�Y
�[���)S�z��[��.�Ǧٛ^��Հj##�h�2�����t+���-��7L�fd�#-��������&�L�Y�:~���Y���e�(�x7��5���"��Z,��4��EwCͭ���/&�*@�*��/<A.o`���5�H�uL�f������2�q��J)mL/[�◐[fhdӞ�'"2����a�顶�������8ҧ�#_�� .���o�l=�����?�<�E���M�̵O�2x��"�����"����{�/y��l�փ�T�[](#7P�w� dA^�G�Vǳ����/�{�#�(,%����	�����8� E�ε��E2*�EJ��?��,U���w@-H�_������`y�њŎ�fR]�0>_i�z7���V5V�amLi�.E]�2�OCk2�����7�}�_�(�/��`�U���AS�H%�9���k �Y����YY�oG�GЈ��a���?��w�#�E�s��%>ly�ʘ�Uu��67o���tj�4j�f(e��I�/~�[9j����Λ�.�X��Cg���RN����gx��m�o�d����|�\侰��Kg]F"�Q��i�"CO@TKћ�jӐ��������e�����(�-K~�R�Ϟ�2w�"�Wә�(��Xy&�~�E-�-<�}��ʟ���?ON`D;����<�j<+���y��Բ>��1ʨt���=B�)w6DL~�4c�ʂ�M��(W[b�%O��H���F
!�t>��s����,����}�9+��أ������xs��=���b�*�VnÇ5?�K��t�V{������Htn�h�>���V�=��zȞ��g$N�I�M��y�z�i{�sW��ނ�,ޣ�t��R�u�_���8K9oe9t<wt�>H�v��$�ƻXUѴE�K����(K G!�|������Fu�>���֋Ga��;~`�����=��}�*��F=��u����QٚU뀼��zɬ��-�ׇ�Y��<��UD��S�@m�R�FC�������4iL�M�1vz�ع%�PN��o3X�������})���Tc�5�zK�Z�2�{��1N��>I^��v8�8�(e*�NL��c�@VW�����	����I�
D�9`j��뺬$_�g�,�RɨݼX?���j� ��W;��}� ��iY��U����p� d1�$���>�a�	 ��@}]G�1>�ڄ����]~*B����ms���k������G~�[4R*P��	׾�� ������sŶ�ʘk�М��������7RuR��D�)�asayX����n��4�er�^�����ۢW��~ś�2�����t-�v?�����hƤw���X�|�T�<p?�G��������ϋH��'�gQ4�:Hx���g��z��DfSW�K���?��K�B2^Z���J��X�^^���p�����%��f|J�0m�e7qo`�\��w����_�r~@mL|�hv1�X��0y �֘-�Z�B��L����h�7����,��AV���
'c��U|Pejq�>)��G����-�X-5F��jG�Q�uh
��ڃ
�HnE�w���,K;�fp�oN�zz�:�-/��Y�k\n�'9�
 J~@.�n�ê�y��谰x����S�̐��y��:'�,���5Ο���(4Լ^G��|F�^G[G�8I��UHs���o�oK�~:DQV���FM����#���F �x���[h&��]�9����߂�^�����8��\�=������	2$�x���:��4�k�,��f!⁉�!y{�X�揋_�[� M�ti散��h^y���B�$|w���V'��pӫ�w�s��ywN�й�*�SkR�l��\�P"4�Ov}��jȔӮX�}��T�r�\�����SY,Q$���Pk�[��:���T��5�f ���|F3�]��"�,�H[�N�O=Tg�n���!���[}��f{��艔J��T���^����5��?���^I���8����#*:�A5ج.:�M�t��v�.����ݽ�~�"�G�w�NȕW�5��0���p�U�־Ky�}�c���ư/3&/s������͗W�Ʋdl�Y�L�:��}�������%�q�H��nR.�:�wc�,~׏S9��ߍ�ϳw]�GZ�Sp'Yy���'�|"���=$+���z�?s�J��	��yo:^�|��l3�v*`���P�I�K��&]\V/��T�����e�`[��ԭ�,b�^��r	�����0h�y6F���\�~F,�#j�I-S�MkW<^(�4����Aē\'M��������
��z�3�B�Ii��q��/5�L|��*u*=�8B@i����teՔ��[��җ��2�x�.���\�|@����e~e10^B�3I�����7���{���������ׯW�f[���*uZꢄz��������ᰉ)N�3,��#���(�Gc�*
1�v)����n��j�1��8O�����ܯ}��O��!��؇��&�����}���}Z���܋�i�G��$>�;��K� ���d�B�����I�eY$7�#���9�xS�[�g���֐f�k;�MS�h)��M�J�m3=���}N`��P<� (�����5���_�
Γ���ꓪZ�5����k�OIpY)��7D�fِ���e��%"�E���l(�_pww����v��6j��uϋ�1f�`��?N3>�^72E����h5;��Z�f7�'q�u��H}�	��I��IW�x�Z�B�ў3*��GC����f$o��e$zG1�56��%��:�����iL��WYѦ���A���Vm�8��[�O\ծ�dq���;,0�Ǩ�k��,ö��ʙ��áIʧ���%�3� :�A��G��=1V���ׯ�R��ς9V�	���|ۓOԦ,0�r�+�j�lk0h*�����F�ܽ�SB_[�t���k(����L�}��Sh��3����DxA���s˹�hV�LI�4����˖���Y&��uϒT��Y�}J�Ϸo�a�������=�*���#�O0�gG��5@����{O��~�O�md^+*����yH�TS�T�b[5�����/J�m��3Ub��q�`j��M;�7u����x����X���2�a���9�����c���	�͇����{$x�ސ�	�H�D,i����2����Ǿ<9�GZ׏���,����'���<����w�~� �7��	�/��
j7?����HN2�(��?��ʉ@
�H_Yr0���&�_9�d�K��TI3��fc�k�~<���f]WFp�=��[���բ}j��ZOP��i�M�v�z�k�՛�/kv�x_�HH�L� h���?hw����
���oln��АrOݣ�'�Th�E\�/cf4�T�A�j�
,�@4����+��R�n��6Ɍ<���}//��(�iOҍ`?�_9�ă`�Ǧ�Y/A�c�7�j%�,�	���uw���py��	S�Kz��cۇ�t͍�`�O��h�c�b�t7SQf��[~IB��;���	�{*W�*`V����OZ̍�6tA�O���<�C�]�=�R��Ӹ���}���8���d�O5ĉJ$YBБ�"�~��$���g_vݬ�j3��I��O���	ރ&x᭖��c�F��đ\7w��\�}p	�ޡ_���PJ��]b�<���U���0��OҰLWL����DdZ��R9��8e��j��+!ƑUO�ln�m�H��6�q+�H.3��1�����Y߉�4���i�Cct����s:v_������2��%�X�y{�����x�0N�_�=P�g{�s��T�݆��m��?���tJy�"�v�U_�+���fG
Xn'��@K^6~��QՎK�ҝU����Y�z-�e�/���%�L����g�WU�d�xsդ!���+ǫӣr�䤌���n�������v+��?�ug�&��eKʓQ&�a I���q�@��M�}<��D���}j}8�ilb�.��L�����]�ׇ����u�^b`�
���'���G�,���j��g���?|���ﶦ�����	��<J ~�q��d7��Jv��
��踿}Jh��\$�������Yc�MH�^��%$g\�QL�Q�z�gT�|���j����ࢦ�Y�����	v�m@�M7MC#��x�;-<�q
���]U/��!S�y�����V�m� ���C�Nxa
G������J�/�|1�^���2m�c�g�|��f�iV�ލ����&��^��2��{�c���d�@��D� =?�[��,A����`�iz��eAǂ�5���󼱟����qw��J�K圄����Ր�{g\M~��<�Kٷ�X�����q�~���y��n�G��F��w_�ee%e����a��l�Y���a%us�nh�ޙ�ܕ1�+'/%��%�ٞB������|��vS?��&n3����+�}P�$;���qCGx������5�/}������A�S����]Q!J��F����X�8���EeC$qf���=��= �pV+��"U��kKs�ʜå�%LH��(~��M��Rw�|��7����^�}}j6L���:&��K�� C)>� 2�+Dq��gj V��C����h��������K�������&FE��:����:t|:7���r�;��s��8��Z7��F�����	\�#���u/VR�g/�?U�'�J�(���>tL3��9!� y���29�	K�Mi����]�����Q�O�����?y���)m��^(��Ћ T'��W"~���f\��y$��++ �@t5���
�h�-�.8꾳h�gA��	!ΌW5��%�\����r�b2c)J�i���t�w���MH���R4~b(i��~�7��W���{��Q�-,��Qx�W�}|887��L��#��E�w���q@`0>)J���V���K��nJ?<���x�Åu�0����N _O�YX�y�ۗ��_�}��, Q��m�������a�3�Ӄ�'_�>�o�����?�
��R���ZC��*��o��z�#�O�)��^J�Xrb�t�UO���rk-N��m�H�-KM�_٭PAm�p݁J�''�	c%$�y=|�Vc~��<��%�)1(L���7���fe7�){���>�-���ԛV�<�� ��%���'�0��ZD8�D{ ~ �|I�u��$�t�o���J���Bw7Ý��2����f\�ᙼDݙo����jw �B��:ǽL�f{�>�Y��l��s��nsO�}k[q��;J��M�}���bS2��)y��8)�R+��j��$�M��-(e�*C�auo;�ڔ\u�A�Gyx�Ѕ����'��2����t�����j�fd0�1eg_�z�>V�u0iKs�/S��+�������7��{��� ��Wns=Ɏj~X��z�D�v��������~/��J���m�i�q0�'���[�л38�Wz�5�^��gH� �J=t���n4�k�0�x��%�F�m�@P��[������Ps�"�Ʉ!tR`cʭ���,N��Y��P)5�-fz�������9��JV��4�}&%�Ɂ�T3��TXt ri��=�m �3�H�&�iI~�d����ή^��7=;t�$�Od��Q��]�w5G���'���D�
}|<��R5釥-Y�N�@k9��}�������M�/��n���cr��c�a��nx��o%yT�n:��Ά�E���9�'������-	7p������U;�>x�C�A%)��9|�����W73�u��s {����7�/���|���`�y�h֫|Ļ��}�W�����K}x���?>g���H�lK/���~A�5^Q�@�g���֧�a�ۀ���]0
hh6%��K-�8��V�50�(9�o�ύ�ƍ�׆	֌ȏ�a>ly�%�x��Š���A�''#蕎.��`�$��U-�Z�Oއ9�~t��%�J����I�5'�u�טVQg��5~����q}_ZJjk��;����
��mg}���	�J�W��i��C�С�����@������)6�a4p~twfs�.���^��������?���5�4�D\o:p��^a@k^�$U7��C�%�qv�
�V[+�1�n��뻩[���n1��~�y�{��gnvn]���6D!w�_����u��k�1�����˪07(�MҳJ�Qh�u��;���H0)�?jq���/��a8��k�&����C��zFD<3W,���ij�}ei���w�e�?ӧ�br�w4t/�DU��L��q��U�#mGD���Y	�����j��[�N0�h��Wb}��t|�
�|�Ed�V(�}�Vy�K�/y�V��J��R#�%g�R��Y����l.���y�.Ǚ��Xк�v=Z���0P� ������e�6f'��&{����������Ex��џ_Պ�O�'P��2��؞`�x�M9A�lv��c�~Ȑ��|�V��7-��z�E��-"V�pD��Z��~�cܔi�/�h2�$݋[H1-�{�bQm� va�B!|ģ����/�4�E��*��
�2s�%<i��f�����|6ͷea�_O����F�4\��3�ȒKN�Hص�e2K�����1%is��5xv@-��~��`oŹ&��d�%S�;451�S���X���`
SR���9�M���H�J%7��]�i�IT��f.+�E8�w��2��R�L�_�\�{ �}���{i��_�VP��z��pFw�Z�Jr�������4�,Qm4��GD�F��z��2i(�UK?�,S\���!6��FT�M���ߒ�};���CD5H0�_-�&� ��O��buy���G�D�{��K|&|��lBgl�Em���
?�Wdp�&��Ѷ�"���Y��f����ֆM=���z�����i	i�8.�G��G,���rij[��m1�ΝgMU'�|.�y�����;fk,���_�Y���	�M%C����2��uP����C� �<<O3��p���΅��p򀫨�"�&��m5���D��#�g& \N�,[v�uI�zA��5�����"G���W�����ؠ��h�K�G
���+����qi����~..H%��=���X���d�|�W��=�5�(Ӆ�3ҭr%t�.���s�Ua�5]}�mY,9f=7z]0S]R�R��@����?�m�W"�vG��u�l"�N��8�S����m[��<|M���W��E��(yn��
7W֥D8��I�NI��+��|�v���<�}�����?��f�_b
�����Cn+����ݹD��nz�v��	/U1��V?��U�A���4l�砓R-�R�s�q?yb��>���.���� s[w�=�Ӻړ]\�̀�x1�_x���l'㾴L�`o��.�G#�j�����@�o����8�W��c9����u�N�l$F�7I�Y��O���s=�����1�Ewv��܆mшa����\���pT�z�wh�R���K��TU�$Lv�<)�k�Q�,!}\��h԰���Q�0�~J%-��'7�É��`q�ΛL�'Vދ�%:��RA�@`�6��Ҩ�\�d�*Y��}z7����ZM����A6�o[7�v��ض���jGJ���Kk�6��T6QTF��ݯ��L��#璘�V����Y�dԕGo���{�y8�K�'����i���!���~����^�|b���v\ǵ�����K��`bnU#�/�pBԾj�Od�$�ٿ|ǥ'��>)���]���x5��m�Y�\9#�ױ�rr2�l�����Q��ш�A��B���f}m���q�
M�Zɚo ����#�Oz'��d���t��
������;-�͝
���ZЀ��/�K���C�m�,��|�L
�P+m��2���ۯ/Zn���A;.�{>z`�\�ED��w;�'���KV��E��a8D�����g��R�Έ�ň�޷��n�2\}�г�r������b=xw����t1���O&�+���dn������~����NF�+���K좇��Q�_�舿%ELGZ�n3B�zn�o�dD�/�9�,7�A�#6��
�-:J�����^.���=�^.nr���Tr"~:s̛�8��	X6.﮺�Jp֑M������V�t�8OT����=��9������n[I�����ͣ~[��#�x�~��b�E��Q�,�p�0�7\��������C	���<?1�=��)�[���!��U�z9X��
�����S�`�Uj�2��h�`�V��OJT�$b��������8^���{B�Ube�h��rgP�$��$�Rd�����lԕ�^Q77���"�݅���e��I)[١�띔!�g)��_���!�������}�]J�lm�S�8��(��*�E�N�A�^��~o�,����{��f�
�<�� ��z��w��/��/T���`{j��Q\o�+q���6Hb޳��S9�[:����.\c|���&���3\�[)9�qE���q+�!�\4j����ܰ��C�Y�V���y��Q�k�
µ�F���:܇�Ӡ�:����s�$}��'�Z��({x]�M<w��7�h�H"=`���^6��ϩufɓ�Ӡ�'�+��+���7���li{�)'g2�=S����Ц,�z����x��;]���%�& ��ȩ�dp�2�Q:����{�&	�x�Xh\��KG�M���3���j�=������-B���׃�����=��7�m�g�w���O�fi���d"���WAc$S=��|ֲ32�G�
�]M�m���~hp/h+�M�{V���a|]�C�qZF�tWh~#ݗ%�8c��Z>�m����<����:��]>�pz��R�z>�|�������]?�܈. >�!A��r2д�Ho�
1Sד���a�S�����>��X<�QJ��I����_�������-ԫa�q�w]S�����{�!� a�h�9tq�W��bǍNӜEa�ت�&w��k���$;�lW�8�1oG��_=��ߕ��o���Ii
?k��� r�
���~Xn�����J�}�J9��.����
F�M6�����>�8=9�sF�W�3��c���K��֐�K[�v�l"�p;�N����M�9E�(�z��A���QО��� ��u��bF5�%B��X�)�~�`���:`�U��X�4wg�O��zϧ�s�9fu��&\��;S����av9I�#�'����#������.�����;q�x|���p�6�s=�o�bS1�G����Ʊ�ZN7mNGG��(��G��헌l͵XW�r�j�v������hv�	���*� 
ڠK��HɹB�c��c�sQ��cT^}2L�k~��|L���,��Us:�a�Ț"C,~��J�<�f��}/�k�i5=�v�9]̀/{�i�w�ϗ��	�@����� K^Y�c������'�/�9���6�R���L*��[y��.���P_�n���sп�&��oq�]o��׺u�s��\?������7p��R�V�\��}����+J�-ɚ6eL簋�B�Lz�x�i�{瓺Ք̝q�r�䛛�	kRN�Wp��_5�c�_���aV���b� %�Kqu�u�J�Ю��_�1W��Q�n��9��.zs��'��
��P*%q�������J�G��P�*r��n����L��S�^No���Ы���@��W�g�4�Y�c׾��T�y����	� ��w���U'%j9��D��+|�7EF��h=�+F��lLI#��(���e9vhחϭ(]Eآ���k���b*	S���T��e�C��ޟ&C���j K���O��(A�bP1�����2���U��=�"r���^o��-�Ih����P?�.��U*��F�H����bF2t]�#�6�� :S�Iu+���s,v��8by�9��
CT�B�E��Q�����t��;s���@�� ����d�!8lg��=}�J��s2j@��q�n�Q�kQ�^�֎8��m���(�������a��SWF�Uk=��f��u��%���3��+��kY��H$��i���g����g���5	ob֫p��l�Hv�w�^�ބ�����3�$ǆ338�&��򆽯`[�Kg�,<��E��8�^;^i7I���Y�}�Ӹb}i���JRT���@U�����қ�R�3SQ��Vo�+��y��:��	��]�s%G�KF3��Vj�ס��o<l�hl�'��l?�d�(	%�Qds����-�|BI�=ƈ;�E$䶃���O���z�D�,y��Э.$���~o����5�����{�����J��"�������LRꮁ���;_U��*Ŷ���j�{پz�.�
���M� _F�����2�����u2����ꐎN3	���A��jf�7�e^�CH����Z��B�
Ɇ�Y�N9N�7[����3�w�X��w��D���)]�>з��KLxLg��V���=��dhByC�P7�P\�\���ۜ���=��p�݈2(�������*!n��ˉ3��t�C^M�;zvB(M��u�J!�2�(���
/�$P�L��v�L���햺���}�׈VAN=;'RLa3�5�7�D�,�p�W�{�h''l�,����`\\��${C�I�,uQכE�������c�1����bb[��Kk��5��I) �xD��{�'�6����"=̔,���e%�?rm�������5�"d��i��}J�@aaҭg`_�S�<�diku���xz\�Ѥ��eP2vc/_~%G��f�L��W��>m&<d!���󡥖�!��-�g��Oc���c�K��1�|.�(�D��Vz�9��
�廦�q��P`�~F |t�%Z�_����V��ϻ�?��0[C0%~��E�X�Z���O������P��!�?Ҳ-�[�����\|k��2��p��)�D������cn�~r*�"��&�@~��㾯߫��ɬ�I�K��e��_�C���|x.�:�v�,�?[7�>^�Ĉ�R�K���D�+��2%��d��^�:��DRy�"
�|P}���%�����-�bn��Z���@�`�](�M���p(��_�й;�t��C,���k�O�����$�X�_2inE��	{��Wv�1�ol�~�RxN-Z��D��%k�9�o�`{u7����w���Q	l(���m��j�z|'X��b���� �E�Ho�(9���:�e�O�CIZ��̏Ԯ(��c��{e�1�����~�2��rR���,k��X@՚���ǁ7��2l�1�O��Z������8� ��r��2����Se���B���4M狭���|)i��U�H]r�/ ȯ'����̫���?�r5$c4ct(�� �������ʠ�5"˦�����4���e<��%ھ!m��2��qG�m�eξ���xi�E���#^���������{�29?�����c�0m47i��O���G$& �a(q�v� �#��z	�� 3W,��,�����Γ�)M����ڛw�%kt���G�g���y>kUf��B����~Ra��\t�����	-e�wa �Y~�_ӥ������bsQ��x��ca_�xhx�4^�O9�@DgBXby@ �9kuo$��y�������V>���s�h-�c$�y�da�Dz��{���6Ǽ 
�)Ru��;��E��n�۴�ѐ;o�""2^WK�&gC=�˯c���~nvZ��h�d��E%s��g��ٝ�4+�҈�ތP���&��c��&b��߅2i~_\>�@^r��Q��9@x��qhx/��s׮5����VޜE��dC������rQQ��#<P���d0�=��y��<mv��V��0	!��9�T�5��~��e� �����2v.����o����m�VKJ� �>�>d��!|i�%\B����8:����4�L¤�`�qY�|�U�&��5
qXԾ7���']W�������m��7��&�%	��YE��y�̕�Og���]`՚��7��K.A0h6�- P5���Wu:�%�.|��l�e���ѭ���'��y(�N�t����I�|y�S�2R<v����w����: 
	��]K����O�Tf	'�����s�Qg�c$�T8暠RM�[����lM�O�鐔+�뎄}�B:�W$�U�ķ:Sh2�)\5��*�},���廓���Ax�H8��	零@H�%���2	�8�����]ɘs��/lD�6G&*���v�I��QuM	9D����W�-����Au �d���<���v��k[hN�]ބ
u�2a���\�H^�T���G���X�KK�6c&�n���\���'��,s��"�D�;l�^ ������K��u[��`S�\�1sϨ<z9�I���h6��z�Z�5�PP̰O��uPx|I�*�Ov��|��+�}/�8��q�o[5!D��b�<0í(.��[r�I8�4x/��Y��񟠐ɣ�Zd��t-]���˘ՔrQP�>�.�o���>m׷K��L����(y d�������u@T�����X���u�?��G��x��ǅ�k�#Y�/9�t��������a«�Ϝw.:`�H����D�`�=��g�j�'H��.�T_]Z���f��"���kps�LY!q�I����Τ�����#畹1��E����l%*FA�.�ǧW'y�殟�P�Z�Uu׹����<��ec�A���x��n�|O�z��X�8��]jՙ�k"몋�g��~L��w-��1?�=�,�;�,����y�g�_&���A%0J������d��\SЛ?��{MJ��M'
j����:Y��6g�UW  ��8_���	��ܜI�@U���D
$;���C�5b��bMv&sʴKl:c��8x/�CPw ��h${�|G?����"l�u����o������#�BN���A�S�E���e�-�!dgO�T�:����	Zl�9@$>�(�0��
D!���ql���Gp�$_�� ��(T4����Bb�E�C:k�H@��v[NVG`� #��Gd�(���o��c���"-�B���튾�z����g���;�s��5��h�Vʍv��d�<��2sD!�eFXÔ��הP�b�Կ�/�:U�L�*�T��#0�o�H���ݠ�iDJ�[�Jl+vO���5w-�T�$ ��e: 57���6?���5��h=Nt�I�7p�W;P���x��EA[�F����%'=$OkS�X�0��v�B���M\2mc��[���<������m1�U&�����H�+1��nt*���J����Q����j����z�mY�ԕ��x�Q���������fѲ�@u�&u�P&Y�°��{���H�6Y�e�Q�Y��!!�Q��z�x)�l4��)���͞�w^�`;�50si�im�<�$ga.��`uQUR�����~"��$��_�']��ݾ;,�N���6{i�r����5��
��%�5����lz���$�&^�^���e��0���tx�2��x���W&����!]����[<F�kI1�U�����.��*r��q��EMA�T�R�� �<7��-xQ�t���`"�Kv���U��)�N�(.`��~��Y��T��u׻��.�Ce���%#dvO���Gqf{H��f#;@|F�WT��	
%���Jv'z�3�x�"De���oR�>��{��b b�tfה����A+H�	;�JY�ΰO�]� ��LU�mHA�H�ؕ�ć>�9�=g��)vr�@��q^UW~��@R��U����\ƲCǠ����t��265)���/������g�3f�>�����Sx�!v��l��𽋞 (��j̏ġ7��o:8� �\�5 �O;+�����w���J@�p��OþON�x��h�Y8B�t���?��U�!oqi�5��Vu@%��J:��A�VP���g�3&�qT(�s���c�"�i^<�?����a␨�zu�vv)�w�m��r�2����Wv��@ Jb~P8L�ŷ�����	��̍T��J}��]Z�_�+{�6L����Sa�ܠC��ki��m�羨�8�(9uRj��j:m]���3-]�ӑv���ͺ��fXn��)�I�̹^�����^��V`?Hj��'��iе�g��WJ�0\o���$��*w�/_ڻ�	O3R�牟|��g���W(Z�P��<e��^�ն�u�
���<�JO�H�~�%���R�����x��_O]�a�**z���
l�q�PC���γ#��)q��B5 ^� ���v��6�^巵��a�'���J�
 Z�'�x��K�����rwG��[�4��7��}�I&���Sވj��-y�1��|7�t�JI����χF���z�����b�"�߯��zPF��<ψ�:��O�%E��	<^v�'B_%�<1�B�O^��	�����g�K�ڑt"H8�\��q?�����~=%:%�`��z����ϡ��E%�������v<~�`�T	���fm��Oc5�I���z��V|�ҧ�^���Aʾ>����}g�+��g�⋀҆���|�g�����g( +Es��k������np<i�l���}��<I�
�nu� �7GI��JX&��I;F��D���sF*b�Ƅ��䮏
�}�z'{A���6(���:/I��ovd�Z��Bsq�֘�/�%������*�@�-5ξ��ċ��|6���d�;A���dd�IWBRmO�1%���v�K�Ho4u��hT�yu���3��`��r���y`gӶ��L�����'*8���O�[T��ۺ�R�
��hܫg��SA�^st�3�4�|-+����X�qԽ�Ҍ}"`�Ϸ��]�E6�4�8{�΃�$��.������
�&Q��=�wz�c�[�����ʢ3��Ы'F�BJ��.n�"`c�Df���r2�Obi�8����0�yL֣�+3A�;=�z�tu��r��@�&��&{,Q��ΨM����w+(^�.��hh�,�DۚD$�P��bp��ty��l�r�t��dq<S�x{9zB�;K��^.*�f0�&���@��� ���ҋT��S��Ɣ�+댝�[�i�WO��,D�Y�>O��J�i��������w�<2�dq�L�{w!���En@H�b�����
]�o��j����J�PR�.�򴺬�]s7��#m�wЪ��]+��	����I�4#�sr��c��32�Q!:B���d��Ʒ�������ˍ	�H�C��jw�a�Po|n˥�nҭiنj���K�|����uuƄkR��!�!��l�:Ґn�.��Mf׶wxQ�.yz���y��Z��=1����U
=�z�#�~1'��\�wW����V��2\}�K5s=� )Xck|G�*L3��moWٕ�ix�?a��P5��	�/��oH��<�l�a�kL�츥+]��F(��j���?���]98X�?#�oD��Y�L�����DrQ�2H�y��,���/����la@6��B�E�����2[��\���>ꎹ��7}x�O�2��A�ʍG�aoў����սL��G�[���'����j���B���s���cV*�|'9u�T���0��e��s��ͥ��x36��Ǣ��W�
�.ɹL$�������y���(�<�>IUp�n�2.W?<,J��~2���w@;���y�v�,M��buC����Y`��o�{�#����-[�o�%(��,m��譜���L<������^=	F��܅����������mav9��bj{�=		���6Z(ՋEE����24Cވ�$9K|�.4n�zua�yl϶��9j������y���Ӯ�ԡ�gR[���T�s�������h [��#/nK���s�uHK��0t��wd�%b�Ou]/,��Ln�2Qޢ%�玗.��#���msmh���v��:Q��-J�S]ؤhl����q~F ��BU"ř���}�ku��@V�kN���u����ޞmq9C��r��uG����t*�S�Q���l��L6!��;����� ����C�V����B�����~�#Ui�����oM`[�=#�̱ ���1�E�qi��t@�#%���QaP����Q!�GG% ����0C	�~���ܿ�>��od��ʻ޵v	�"�zV��FewR��h�|����]������l�v��}h��S��N��N�}! ��+Ӡ�&�y��ǭ�t�~Oi�a��3Bҝ[\�K	���a߿���������"���Vg�j9��/I{�+�s����/��O�5L7p�Y����g�9��m�������ӝ��ޜ�#�H	i�$�46W�������wt�\���/I'QFF2
Z�M�p�֐������g����p']ϓ�^]y=�lc|7�ǥ ��ش����~�Ѝ#���,���F���*ճl��1����՟hY x��};���q�N~X�<\��T<�t�a�)9*���f$��{�CR>���sq?�ɳSV��\1��-�ҙwa��V͹aFh}���������P��yqR>H��6pW�O�|׍�0(�> ]ڄ�"�����A�u�n?�ߩְ�ʼ#�t#Ь�)Tf�	�x���+�g#�sV���x0��Cr`�"�&��'V6��cg
�.3��o�A4��� A6��.��'o1�Lذ�⊭~۱ޑe����;��
�5�����'��VHhQ�Ph�>Zl��q0� I(�la�B�G�o
�*;xtwoL��1@�1��^t�l ����*��
`Q�� ;Z��?G��EF�\��m]�+9�2��o1n>��H'b��/g٘+ndn1�9:\]�[���񤤰}�VxKNI�K��w� (��uC��-�Z��@j:x�񈮼�1Yk{jgs�mip ��/%�w9�[#ۮ�f����a�& ��駚�����2?�Z'_��|8�)Y� �����P,���t@JhrW��A�7!b�
���o3]�������ʺ7>����^|I�[�v�����n�6~Ǒr�7=݇�2�?@�����#���m�{��
���j�I���p|_@%]�:T6� ������K�Ev�A��+�y����U���y;�hZ9� �0d���~3U>G����"�
�5Hm�%�F��������G�����ĔU
��4j�mo֐��2�`?'����	�i�\���3�bUS=�K_�}�
m	o}��@����O�h��`�ʦ\�����L
�&�����#������������"�[�_@��Ji�&'�}���)�x����?�01W�r�4��O6HS�6�c���|�^�o�9�!�X�T�@�!�!��� ��M�V[�j�'h20E�N�*:c.�᱉eJb�~��yހ?1�)������u�2��.���34c�aÃ����n��9��g�Zmo��� �{+lO�ģ����&�ʁ���i/��'��q�*AYR_֟;�c(�D's��C�x$�M�4(��h���6Yk[8��
U���^�F��`���a������l�BW�/ut��M����̛<�?q�*���Je��ﴞ��!A����]�q(%	� �%%�R�I�ہ�&�4�������}Ru���9rG��|�KIA	G�zk^�A���$f(k	A��gx�W�� �����ZSۚWLr=@b������ �퍓ɂ�jI�?)��>��_�w�1ĬF�h��Auhn��a����\(%�	hvK��v$��@3�+u=��.(i.�;�b�>���UQK�:R^d���o�ȁ,�f�i7p0��c�x��`K+�kO�>v���j�
�Uɸ�t}���_��R�D}GA-
FWo
�
�1^ �ڟ>"lQ���������4jr�UT#x8��8J�-Zp�xv@m�_W@���)����-�̜A�æ�ӱ0jw��9�bW��`��Eࣀ<*�W��-ț���w ߗ���=}J I����;��y�e�}��f���ap� p
�6�!��lO�⏧���C��H��)���X�Q`_m��_��+���6�w/M]0J��`EΙ�Ԛ�`�l��;��g�A�\�f�9/�����Zh���)�W�7���رƈ�7vp�M����,K� �����] "R��?�������^rV�T�F���"�{A/�:(����\���	��Ȧ�N#{�N~�X|E�yʦBi��E1���f7jy�����O3���G��y�YV?�66�O2sO
�����-�H�c��!u��B��V�=�5+�6�ݘY�W�����c�Xv�&*�A�v��U.r���폚]�7Lpo�i����k�mڳͳ�)#ߢszv�j�� ;��HҀkYpc�|J�w�G]$[?b*�o���"_:���Xۡ�9�1�7��-o�����	��k��<E8�E�#�O�}��������+�Шm�r	��Ja�e�I�ԶYmYZ�4��R��)��B���^ZB��t��4��ݔ^�)�$`O9���#j�㖛��N�E;3~Vhw�+ħj�y����r�ޭ.��j��2�������O��C؂�IU�jo��fVH�l����OqLo���tр�ᨣ'�d��#
ծb�P��������++'�7q?
{E1�h}]� �#>�G�Q�=���+{BTM�zK%���jӋ�qڍ7���	�>|�
���4@d���
p=�l}�j_�Hm�˛;�R�z���RÞ$WS�E�@	�G�b;�j�s�o���5A�,��V���4��˔#�?t��l�@)�Pk�:t�Ӑ9�-�[(�'Wa��q������{Q+��.�����Z�Ŧ������(-i���[<��IQ@��iT7�h���Zv��3?
L����y�8�#G�L�쉩�
���2��A��y��#�̋s�b�`��^������	��r����ڨn91��]�i�8W���l,�>An�,��8t�\�]�Q��'!D�C��a��Q�.bl��kLO	�)-�S^P�WnEXD���t�mw�H������r�i(a��:K}���R�)*�T
;�J���%Wc��HDy9�.���H#�l�N~���ԍ�W����-��[��R��9VD�����>5f��`W�G%�|{Brr�\�S�"%f)bm:#���(旿y�t��wMsB�}H�ǖ��+lQ'���ز���7�\�	=�V�	����vͪ���Q��l��c����J7>$n����0B���nbF�Tj�a;�iޛ�cիGKo�b�־ƺS��������H㦨a����n��u���_m�k�<�j.�1xi�d��O�o}T�b~�B}e�L���DG����P��]zQ7mb�t���6o��2.���?�4S[�<cɅ\�G�����o��_�a��Dr_QvC+]Gu�3�}K #�\��Ʌxëo��q���Z6h�gr0��ϽԨ��3�{7�\��lsh��0�4�y�;�VN���@������P�7V���N��kf�fpc��p�rխ�K�����D��oR�,f����d��;'}��гue��Q�a`�b�������x�`���^U-1~�ϰ�Ϳ�]W��Q�j��kO/.�};4(8�j�0�]��(��y��'[]���y��|�m���I2h.���	?�B��/,0�t˸�$3���O�~�)�63�W�S�i�a�'�&Ҋ���we�MJg���ʩKT�<W1Z����W΃j''�gf�M~���rz8̞hg�c/��.V�����y`�c�7Cmߢ�|Æ����V����P.Q5�K�:������I�:�
3��q��۠g
���J��Tcr�z��*��Q����baK�,<l=����鄟��a<�q����k�i���ư�W��T	����@�$��4$��. ��N%�s��$w�#��4�3��7r����đ�d��p�
�gF.�%�p�D8��b��%uz�b��d�G䄚��`-~�=%�ɪ��~�u��Ah<SF���On�B)2��%�7��g�Î�@0�Vr��o$94dbw=3	W�ݤ@�%���ri�)�c��:�XI�w�����=��q����J�ѺW!X���IYY�ۂ�\�Ny9�t��)8-#>�G��:Vnm6/�{�J̛�|�D'�CUjR��;�����aL�a�q�ϫ�ʲ늱"�BIFi)����*��F�Gӌy���S���,o
B�w������%mKS3yRBڟ�v�^T�v��T-&E�V<.cf̭�u�bw���T��x+���"�d�*%�i�ﾓ)� �<b��x�ՙ0-%����tfTcFv�X���Џ$tx�Ҡ��&�ha������Č3	� rc�ٍXL�B�*�Ж^?�G>~^��������(������P�O
r$�M�?oa� Z�)i���������$OPޒ��(#�;!I�P�9M��Y�/���B���'��N�^zq�S!=_J��߲o]5d5�h���U�3:Vݵ��<c�Tۛ�,��S��0IZD������xl� �j�^G��{�PW[��\r�Qn�%��O~V��*4A�d����2J�#f$xv�,E-դb�#�5|rD�'ޠx��n��>�b)���NT�p1Z��B\���')׎D/�k85v/�?l�Zr�����&�,��KJ	��֭D+�ː;���$�骐s6X�l�2:�s�N�Va�!�W\LD �U�{��7 +��aY�P!��gH�(��3��B�}���XIfaw�T�3�+73���cBe��UЅ��͵���f gj�Pb�_ס�%
��v�h�1�O�37���r��YU�7��O��	�MQ;"Ͼ�N������_��*��pT��{�n���9t�8)�4��%��n����~+-�h���`���g^hD$�(+�^g�j��7��8�J	�y�F:4����ʠ*�uKq�j���Pp�k!�!��x&+"zג���K>d�U�h��~��#6��<;��`F4��Y+��G��%�.�9��M�PK�s��ߍ��d�'���֡.cH^yk}�����T�9�IVr�{��y$��k/eH �]��.��
��pEe�	�k���q2��sB�꼚p�H�ctONg��DF�>�P�]�q�QG��z���BE�!�	��]�İ�>%K����K��H�J�x�憚58��x��W���H�R�@��	ڦ���|����#�͂�=��?���5�$a��fV��@�	��մ'���kk���'��z���dL
y9�p��N2`�b��0X7Lu �ȱBzӵT=p����@ّ�P�&ߩ� ����ޞ�k��M7��8��F��BM4���6�X��y�Tz�4~ܾ:��F�>�	a:c�۝�a�o�>,@��'1�h-^}�h����z��&�$p���=�Dޛ*���%�]Q�b�C7e�0*6ϯgE�����P	���V(����0�=��M3�DP����k�T`�/)�Z�J�(e�������Fr������W��Z��p�q��0�y��ʯUv��se״���V��ई���Խ�!�g��e4s-�\�����4z�K�qU��s��aĭ��ˢK1>TǛt�i�'��kLҰ{Q����iLr/��9�o�����Z�A�|U��~��|8=�[O/�C�J�r=}�����qMJ����z-V u5@��U��FF5��F�Y�F�bL@�LX=��kl�ə�s�	�о��|�`�����t����pB~�%�J�Bkw��选n�U���d݉2����b���ѐ'ʸ6C!v$���k���SSח������T�N�>m�:�f��T���K�:���+p�Ľ�ļg|�R)��������V�ժ���՜�ݡ��?��[�CTz�a��Q�KYҳn/�2LY����w��R��B��
?�#K����֞ľN
��$3�:}6�}��;����?<-h����[ jQ��v�OR�k��G�����$/���|�ӈ���ѹ���&M���|��{7�T,���Ҕ�'��=~��ݹ��*�S}L6��Bӵr�/��$'9r�.SEH7��G��ń��/%h��	���xч؉�y,�&��0�Vr/s��Wd˻�n�pi�S����\�"K/*��p��1�� E��z������C�B~;�B�Իs�N�H��T���>i�]?�c�Z�a69]����Q6�M��:f`�Ϝ?���A{G����E���|�����W6��MZ7p�"�f/�i�`n!�'w�h�>�g�I�R�I��A]�d9g���欉��Q.��|���4�:��`�R�����Z�T��<�(�/���S���4����K�JHF����^N1Q��5�.ũ�*�����[+�ֳ-*�!+�6&2���ˋ�-j��}ЬXFc��ఁ�β�Ɂ��_�����a/�H�N�c2B�Q��	'S���}�����I�=m�V�w������ڠ��_��6T�����q��S��3p`���^`�L}�+Hd>��Z��B��Z��AD>��Od����ηxm�M�\��$lO�m�K����F�F��h��7J�u�90�l�*C�9��+�J�����=0tN�)6���6��Cp���#n�ژ��{TB�/*�"��x��y���e��.�YWr�Xⳙs��aqȺU�dE�T*��!/N����lav���� �[�����g����Ճz�m#?� Q<+������L�JpwY�ꠉ���w�(�r�k]7*�Vꞛȹ{��iቆFl���W�$͹xx���������:<�VJ�=�}���ӟۤ���{�R��a@:��OcCG��y����	�3d4�S��\O�/Q=����a�y�|҄�|�0/Flm�k=�Zz$���0|���d��f~
3y��E�C�b㓅ir���n�uĘ�R6����o#�����ǧ���dv�EXB�qH�{u����CGӑ쵈#��~��NL�'���w��9꽐u�܊^#q�S��J�,(�b�T��������&�L]���W�N�t�N���-8��+7	׿`��+y�w��>#X�&�?7�X��(�m�GY!C��z0A���+x�~������8�'[:BV��u�<�t����v��F��-�'����-������y�4�R�z����8���-!Z��I߾�?'3RFV�CU�ӊejQ9|	���
�C�7q�r��a�Wߣ}�k١<�ƃpMu���%ևu��͏~���y�ԫ�����`�����U����
��Q��I5��@;��"���d?�m�z 1��&
Y��w��� t���d�e�IɎ�&��"��'��m���w�2+܆�.#"���@��5��#�!�gf�aiʻ��0��ޮ�߉�����]8��)��׆LF;�̩Ӭ,Z#�����{��g]�����{��8J��-�����δ�(^y�A�8�?�j�^����	��>5�)ړ- �lp��>�wv[�����x�8%B�s�O��6R#�s�;�͘{�ZS�<�HqpБ���to{s���`�Od�t���(��P� ]Uq]���+�^�̖����_�|S�x+�)>Qx�K#2^,:��=�� |y�0��K�ׄ��'��kC�����Ҋt���x�ʘ��͈G����wa^t���[�1��N�d���!�CR���]�����Cq8�;֟$��X��d�QE���(������
���lzn�.��Q)�~�5_;��R�E�57��ӑ+Vl(�C:��������Q���W�-�XTu��SF�$f|D�ch�/[RyJ�.]�����z�G7��u�-A}T�"�H|����+����ۧ��:���ď��t��#M�
��5Ecs#vrP6=a�6�E.Q�!X��c��1���pHM-	�ĶsD�M�:uN���L��������,w�K���k��[�z=b��~#�;r��e���t�δ�5|ڣlT+��<����h0��T�.�-rԳ@yՈ�F�6���z��	Õ䄿�o��]:�L�q^��Hk�s�k/�����'�Wk��q���KGk{���6��=܉�/7����Z�ӝ�PK   �M�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �M�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   N�X���  �  /   images/dffc241e-8a0d-4217-bd54-7504444465dd.png��PNG

   IHDR   d   �   6ke   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]x�U�~g&�$@
	�PBK I(A��t,��
���eU,�k[uw�u�W*�`�w�7C �@%��:��=��If&3I0�0�9>W��/����v����°��������2�0܅����Ý��W_Ƴ,f9��2�\<tqdbY²��,K4��Ύv�K,ϳ�X}�&��,sY�࡚�؅),+�>�'4O��G��dy�I߱Le����,�X�8����Q�Ph���= "R/���za�7�&Z~P��PU$��/�O�,������|`�n�t�������� R-/��zb�_�h�o2�~�>��I�Fk�
:UG�y��fr�ZeH������������Pu���7`x�������,�X�����2�Fk0|X��CՑp�5�rfVQkl$ChKW��k��0�|��mB/�\UGb�byQ���=/�Yް�#GnohA�tV��ʸ����Ք�͵��I�g�H��,=���Y`(�l&{��qh����@x�b���Y��y,�� U�t�g�3ՎD=�Ƀ^�[�7# nF@܌<��y q3� �f�������7#瀔�	�t:�S�%��x�ܭ�}�&:��[P����{�2 찏��;�Fx��0��� jBޜ`I�9�hD��Mɩ�*�ʒb,+�&=�E��c�݌<�8��ؙ:R{Nѫ�~���I�P�T�p3_� �����+(Ҍz5�x���+�1��(�'/FX�M7VO����(6��Fp����6��:�X��C�����I�p��w9(�a��%�vwf\sU�L g�ƺ��GydLB�����">ə�УM\ѱm�'��}�;�O�X�7�SPPT���uf��q'��D]�c���E��;�C�Q��JƱS�x���=��|��4�8~|�������0w�N|�i��v�㡑�0�G��yS����_�̡��|���۱`�/HN9B�Q�ƽ�Y�x���N���"�ܟ��w�̒���i`�;v0-�36=�F(�U$A^>g�ZJ%/)���	)U��Y�/��_v�#�Y0���IC��F���3�ߦ��f�$M������{Y���䣘ԯ|}*���`?�/��8{�pV�m4lR�#��Y��4@8a���'��:"�K��Â��`�z���a��=1aP?�3zgdb����z�O�=\I�aC�g�!>=�"+��cF�Î�hlLJU���vG����*�}�֝�.��+~BN^>ڶíW�t�2�0Z�)-E�L,��:_P��o�I��R�������2v{j�b�=��p�>1jn��]-�D5���^&C϶-���k�s.-�()v�DP�b�2�M���'���bad�K���c�>��	��w�bϷj@8K(!h̼�p{U$jL�ӎ�V�)��e�R2�)�c�#���
�ye��e�@����]�'S�⮡m�@[��������@t8I���Y�:8F:����&�eF�)���M��#��=�R��+	¯8�}J}N8�ıw8-�\MU��J�v:�͂��>��C����1p��uz�&]���`X�Y�&x���x|��ŷVM�^�������NoU/s�q�sШx5Brf6;�v�A�1���۝M���wmB��*5�rB�&N{�c<��Wj�j#ߝ+(����ց�U�TAI	^]�	[�������0u`o>Z��xӞm=|�^�&�� ���Sc�Ftxh�c:���cCU�lI�����X%Ns��*A��U�d���g���Թ=��~�:�N��J1o�.�QB�5��9��[����֮r��S1��UHI:��h󙰈p<7e"�����\5���4`��Y�疟�BAqI��Oݐ�I���ʃ2�+}�5s8Ƙvm��iHL;�َJ���M�P4�kD��̓z�!d��H��k�H����]	�9��Hڽc�ګ�jH���パ1ј�a�Ũf�5Pb�Q�%q�[��1�0Z���$/��j�H˾�0B'�$&�ge*���Q*R���ܵ|�u�_J�1�O�2�)Y�ۺz����<=�8��9�w��S*l#�mk�|�-��w�Pk��@(/ˮ�R3(�l�~H}�P��Ġ�v�m����Lp�[���`�XѠ�DS�z�O�_ޘ���^#u�7�5hA�t�Hʥ8!=q���wy�h�c��]6��z��u�PŃ�.]�y��\�H]�#h䣂�'Q����z'%��j���S�ơ�Ұ�g�'�*�Y�u�P|�����8K�����+�1�Ǖ�3.�IH�������Jߊ�[Du!�@�i1�ըH������F���SD��hI�����w܌����]/�)z�NL�C��������b{-;ԕ�ď�F}2mI\dD�� ����Lݸ��N�-\	H�em@љ�.��.�����6a��җ�U��6���c�"���
�q�]�lMo��~H��35�ڬmp��W������!��wf�ۊ���(=����6�����9,A�$����^�ڹ!M���b���qXv	e���O�F�
s�����:��M)�e��e&%��P�y7��V"[��*u��+AaRF�����	'��dZ�JM���s`ſ���/f���])G0}֧�Τy24.YgsQ ����ju�\l'!"]Z�i����| �i2��>0�n��Sg5O��w�W���ű$�C��3���hᗄ$�B����>ؼ?�چ��jw/�h� 2����5��/�1P�94��P�6Dd���}Վ�,9��ضK�%��s�t�(}$Rh-�Wm��w}��l�O��NWoųӽ3�w뤼,C=yY"����o��R�]�eY������:8�c!�p��� �Ux�3O�+��6���)uA��0�&���d{M�9 �xة�:�h����R� v��o.��Q|}0�[T�hU&ǀș�.ڠ�����f��¸�n�P��C	�%8�O�D=T��Ԩ�����0���B�_�{��(�InG�W�dn�2��s�2�.��#DpCL��X��߼e���7%�������1����Z���4����C"�	�?76�(@~�������7# nF@܌<��y q3� �f����) ��S;r�qU��L��=һ�.��z��7�܅��*,-�KK֫�jS�؟*'�uq�W�C	�s��j������ ���!���r3� �f��ͨa"�:[V��.G�$i��ʫk��5n���X:&-�����>s���r�=��\xh3�2�J��)�hl��R�%�aB&�m��~z|��p�X���7�a9��䭯&x��)X�;�S)�������Kr�H����_o�9+�a��_��<3�F�0�/I�J�7�R��E0~�'_,R��n܂ןx a������x�A���rDn=����--Ųm�1�W��%r����;�#΍M��E�2"�`�x]�4H@J��%��G�ޫҹ�Y��� ,ٺ��.P%mK<���,~�_Il�p���;�!�"�n����H?uZ1�� �	Bc�F�v���$@ٕ9?��Сk��f-�/-���$ &����� 3�_�+/�2�JҘbԭ���g �}$�z�n�Q_|�jr��{$�eDF�;n�n$v}����pǫ3�G#��T����"-;a���]dy=�D��s�Ԕ& �2�t����	�_~G��{z�x��a�P"ʳ2P�����tu�zc
r�0��>�۟��|��*�I��� 1�[
a|����PDճeO<b���;b}�����G�SG\�O���LA���hD������ �"%͒�&zP���e���%$6�=��X�/��Gye�lڂ��y�dϤA"I�۷�,j�j	Z����X"9J,)1h�;0���t�����x�o�����z�.�v�{b��K�:�U�IRZ�q��<7o��ѮU�eW��W�ñ��xU�uj�޴��� ���ٹ_�&��kC-Z֦�N�} !�t��*Gչ��A��"��J�a�0m���=g�:���(ϭK����?+��1'�����Ø��[�U�a#zw����<R�� �O��=�hw��P(v��u�O��q9c�G'�QI�l�^��*'�Ty�L�l�\و#�(���V3Yޔ�}0���/'~�غ�ϛ?������:�3���v�Txe1����n�A����Od�R׽�x�!�|�I��?�I�������n��#H<z�b�j����LRK墂|}�^�F��t[�Ȭ�Y�2���9P1����c|F�	 *�U���RR��V����=�).�R��4
��?�$�	���9��rx�6H�[Z��Lv��N⃅��ѿW�����T����K����M�۸+w�٬����Y��d���#��/TxZ�LQ��&+5�6˩���m�=�l�eI���ڥ�t������O>�~����a��L���djD�`�>�"��x�%��()�jSIU�93T�+�id�P�Q$w�RzS3�>���{\��ݥ6�Μ�Wu�mxj�|[�.�ը;PU~�����I?#BC��/6e{}��%Kv�D�zK��K;(+��_zG]�h�!�b�&�r����	cɼ��#	�����a����Q7�	hr+�F�Y[X�2��Ոn�Ryf�D�z��Y�@�!���m�wE?�|�i�Ԍ}��5
ٌ�74�urAA%\ڨ������{���ld	��Ĩn?�b`�򗋱���|��������k6!2<L��<J��XR�ۤ��cӎ}���N�h���<�.j�AR�Y@��:��0�����/�2<y�8�eYrQ���_r���d2�����EK��R[aC�;�&�r7�ڔ���I�%��nq�S@��F
D�e��g�#Q%�j�� �Z����G��i�%6��)>>��7+�%ϋ���z�,�X���A�]qyt��R̘��v������n1]pu�nh�;�P�h��;�e���|��^��O��$m�f^�|᳅ؾ7A�Ll�L�j�� d¸!�������%�3DI���^�fR�N��������eر����:9_\^'�:�K�f�g]{����F��TT��gO�]۶�z�+3�G�H��j&W8	W����]�ĝ�I����F�Jj��4�T97^}%@g�lzq��d��� '��	I� ��	��{wǢ����L۸Ǝ��R�Vz$����1J�/e�l�;W��_xB]��)c��T3��yIf|RnB��Z�6��_`��,K��t��Q�����Ć��0ȝU��S��}�W?��D�*<-���V:����~�r=ZRJo?�vg��*��n�c(A�r �����n�7����smZ�Q��,S��5�V��ȭ4��t���V��$���P��������Tv�9�|�LOH��(�)��(�P���A�+�7�]Vyf��M����{��6��`/�ސ�yI�)�$���!�@����.�?]siJ�,��T�I)�C��i�aq�	�n|�h)�fLS��g��#�S�ug��^�d�2�}�:U-=�Z�`�ߦ2�"���o\�ڟ(��!����'�u&W}'��:�kM�-9�8(��=l����"��@X��+�ڄ�V��ȼ$�N��D�֣[g���Sٕ�r_�5qb}A�C�zZ�����x��=�����g����x�QU�< �;D�;e󭯜�Lj�"����gaL�89��8�F9�+�e� �
�Pr�!p��`��z̆��lݦ2�;ї�c g��/6ɏ���R��c�y�*�Qp�!��Y��Z�B`�7Qw>��
�Ibs�4��ek+&�\�$�^n�qb۵US*����;@�n���>[�#�_���cY��Ȅ1xq�oGT��١�1��t2r]Fu�M�E�3�� >d޸�}��#�(�����]2i�@�8�5W��ŝ#����`r�d��x:�b�����/��[�߮ 1�3>��Ҏ�0V�'Y��Y�����@��P6�Is-5�L@�_=��:���&[J��Dn�b��@ �,Yڣ�Dƈ���j�����ӓx��;a��Z~+��a�� δ&�W��F�|��>��v�P2ZӐ� ��vѲi��q%60����:5O3��g�g{&�^��ulO�E^�`�{�n���p��W�>�?�	%jk���jɤ+m�=c�1����iq�%o||�q���W~�n�����b�GYR�����?Q�w'��N�Բ��xq���J��xzΗ�{�0���|6_�e���:n`�؛�&�A�L��٨�a��QBw���)y�38L�j��Xcߑ�����k���o�	ǋ��Dؙ4�p`G�_w��b��T�/�_��R�u?�w����HQ�����^���.ao�N�|��E��MTGd�z���.O\/��͡�V��C�_�7�!�}	a���)_��Vn�^����|n�)J ��d�xwҡJK1��=���v�*��������)�ɻ_o�O}�~zK�{�Jb!�M�j���a$�6��^��;l��r�E�&�>��L��v�YY���e�^���K>������b�S��G�J�����ʭFT��S�~Z��g��񮹄�	�Y���,�h����ބ1��!���>��k��Iz�r�X��7�s�s����8#cFeJ��e�\��I��E��l�*p�gNu ��Y��x	ۧ�d��A�5� q@��4/�I��9(-QI7
����-&�P��,g���5?[V�Ǝ^��U�մ�j�7iEE�� ��mc�Tu���8�(-D��bC4�����H��?� �u2�#R�1�MoDZN+l?_�\�u�}�ք͉}���v�i���W� �g�aSR2A��;����J�aOj7�j��&�qU��Neb����CAI#�܏��ǜ��PF{�=��0����n�?4O�&��8$�@��2 5$�Dd�k�����*���M��51 j'=(� � ��PV$e���P����� �]�����xge�zF& ���q�t֓v�v����) ��ad�����Ɯ��u:��s��s�+�r1���Y�m��^A`.����>�)pj��w]GW������6!�U?o��k{��Gk��O!��f2�Gf�8��8���9=���0���&B���an?�u"�I��*���w1��l��FېU��}X��V���Aܱ���2�E6��#�e0K,.�;rG�8n&�q��|�#��	<��j4h58�$��!M7K}R���t��/ NI��뜶��8#�u:�7Uj����:�U��yP6��DԮ��J&����p�)�р���N[M��;\#��2�� q}�%5��bL^z�'�ƨg�ڻr鴆�̎���	�ر?��U��/v&Q�@dy.Etvj�koRn0dp8CE0��?,�DDW���    IEND�B`�PK   �M�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   N�XrP�	       jsons/user_defined.json�[o�6�����l�i�Ｘ-4�i6`
������4��G�Nb���t���lJ|�O���|�4�+L����W!sUJ��[Y�J����	2-u�u�������?�l���U�U�}9>1r��+]ݛ�#�+�u�T�(d\��@�M�iΊZ�e~��,���8!�)�A��$#�%cJ�KsY�J��u�/���9�"�� ��)�� 	E�XF�SrOV���d���a�n�i[jsc���2���!(��\ի����rM'�y��L���h�q=Jm�nZ�Qy(M�L83���V]�G�0-��p�`wCճ�_��t	�M՚�)X&���Y|���a,��t��'���ه�N,����Lֲqb�����dB.�TjSc/j�f�63�b~:vOVdC���-(�^���&6{Ag��Lm�C���]����_�ϰj�
�U�������_�Ϩj
���,tCm=�)c�S��೛:�(艝���M!?�l��lY!���'Vd?��).[[��b�B��V�u�lZ�/ֽ���M+�Ħn����xR7��X�j�Pc7��F���M�%�o>T�*��-�Iu/�x`㢞T�����zR��"{W�Iu��l^�'�h�?ƞ������a���2G���G$�	��'!�$9�H���{�c� $��W�^ɪQ���:Qs�^{���l+��Q�,a��y�fs���w'�^��3�ą�UV��J޴}���WDV�9�M[c�zm���f��KY6O~
�Q\�+�Y��6/��Y|�_�~:w͕��4�W��OV�y�g�h���f0��@��L�L�P�%q�a�k��3n�Hgf�c�J�L��gy�����qM��ژ��U���)���e� >�V�ˀ<MY#�7�L�.tkX��5z$�j�ؙJgy<��h�e��|oU�ҍ�,����X�������;m��:c��U��Ré������NC���;/�ވ�F��
��[��u�,�����V"����F��n_2��k΢H ���MMS!��n��	5;��lS��z~���������Q��ѧ���H�����}X6�*e3����ڔ~�W�Pf�d0�s� )H0�#�0��W�dI�pC�9��E��ss��	��|�kg:�4��U�>x"<A)]���}��4��%d�	������@�|������7�u�O���/�n�m,�>�ś�z��;��2�_	q�'�m9㷆x�'�d��|�g�s���٨v���SdV�� ��+E�+
������_PK
   N�Xf_��|  �h                   cirkitFile.jsonPK
   �M�X����7  �  /             �  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   N�X���a� �] /             -  images/43b8fa2f-aa16-4fa0-a6a4-ecf006c83c4c.pngPK
   �M�X�&�}[  y`  /             ۾ images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   �M�X$7h�!  �!  /             � images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   N�X���  �  /             �< images/dffc241e-8a0d-4217-bd54-7504444465dd.pngPK
   �M�XP��/�  ǽ  /             3[ images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   N�XrP�	                 � jsons/user_defined.jsonPK      �  �   