PK   d��X�kƏ�  ��     cirkitFile.json�]�s�F��WT�/wUw�}�8�^�ֱk]�|�\*</ɅH;^�����7@64CI���J$LOOc��=ݍ��ˠJ?��m>���GW=�g��5���]Z��ݫd8�������oU:�\�'��s����lꦋ۴4F��Y�Ayb����E!˭��-\��0|tw֝�u�a�to�L*�,�`baI2���RRf\��(}+�皤�2I!�`�Aߜ&��"��0k�}%wJ 6̂��&W*1\hedJ�ߪ��IEYf2�E�'�(hbK-���KG`X����%�&[�L��l0ٔ�6�m6ۦc�Q3hPBR�E��&���󐙧"P�@�*� �i�Q�6�6dh24T��*��Y�.�2�&h�e��6h�@]c���L`��m���w�e���Gu�[吻L;l�\��]ʊt!F��Ud��>2ҝ
��@!��gv�uF��n��y���FI�)�h]d�(�NRƲ$#�ж�DAӠ��K�P���[YQ����a���<p?��Z�Jb:���[`��]�$ˍ��󄛜�J�,1*�)yʴf������dd	�Čܽ�#�� �Y��]�5�O�A��s��hf��(�wE�H��֬cd����#]�2�]�'�եȜ��	2�u�@����"C����#C��!Cw�����w-T���]0eH�,�C��yؒ�&�*�a��?H��n���\"paQ��(\��R��\dYT.:
�8�g&�����H���^���o��0q���`�4�ib�R�!ljS�R,�Y$�,�f�.u�M�8(f&�8���A1?�bl.<�8��U(l������uG�E��9�Ӟ6�A��k���F�r������x��R#��q'IH��YO��pGg-86yyzW��!#p9�KcӃ��s�Ŧ�N˂M��/6%vv��֙;B��"p��|hl����#E����6����&���<,҅��L�rQ���lO8���ED�"�pQQ��(\L.6�"�7zi��8��q L� �Ɓ0��a�4�Y�H68�Y�8(fqP�⠘�A1��b�<��Y��=�\��rV��ٞp.g�	��9���	�rv��ٞ�\�ٞp.����	�ru�lO8���f{¹����lO8�����9m�ٞp.gU ��	�r^l�'�KYΚt�'��YӀ���s9k�ٞp.�+�u���XU�܎�?ה�ƕ{��O������*\5�~�Vt�\�����!Ņ!L���H#���gz�{F�P��i����n���x�##���c䋿�҉nd�O;d�����sh1{t�F�1]���-������ij�����a����;n�2Q�!OiB�1���Ç�sZ���G�N�i�樾!��[�� �i=)�S������ �w���ϻ��K�u.� x�K.ҵ!��i����?)�S��'x
��� O���c 0�@`,p1C�	.f����%x� !|
B�pE�%�NK��C�sC�("���x��r��=[W����-��,}�������	�������!�cqB_q���u�&��1l�h�+�k]�x0�!���
�l]�� ���D�V6��pm�%�AF2�ʆ��Y�bh=�#~A~G(�Y(��� �敇┟�)�p1���'�]��3��zE�7�.\<���c+q���1�t=w���d���	�۵�]ȫ�Ǹ�����1d�[��l�	C��{<�c'D@����8�A�Dp�xr����]$��]-�>�l\t�$neх�z�.�<���kG�R��G�0:�rʎ��BJ2���/�ܲ>��|>	���C�<�<&�z��m���ޯ�7E޺ծA�QOJ=-���SSON=}�?���=X���`��=���|�{0߃��������[|`��1��N�s��� ��+t����@���``�7j)�%�	�
	]M�ӄ#re3�[hX��rY$9,_"�����y�K�'2_Q���.�EN�����te�`a�˅�YsH"I��&�X�� 8QI�gYAt�aBJ��R��9W2�5IF�MT���Xk����T�İF'���F�h�
a,_�AiX�D��9�Tg"q������2��1IAN�7k2���$����]^�Tx�^�o�~�O�<�C�@ �\�x��E�'x���U�kA�����gA'��U���AǠ�xa��ǞJ�����؃�fP`��{v(rX�q��e�����:�C�u�ǉ��o����� �>w�${�,�[\�4s�,�w~v�+�-�i��M�ib�M�i��M�i�M�i��M�iR�M�i��M�i2�M�i�GMt=�x:�f:������6�\Zd�������v2~X�����J>|�.�_�������]��:��O����à�j<�����o�:|L'K��_�9򓳜�a���p7��f�
���t����U�����m�U��q� �XTK7u�N�e�/���N	�K�#ɪL"�$�����xQ���Rj��6�{������ L-2)O��$т�IJ`����h���`�L�/���z/�i�b�
���Y5.�J��r�y��|�e}��ɡ0���m�;����&���\�;���u������n��u�s]n�K��wFȈL�{ELg��Ż{��^�����e;{i��|�Φz�ۛ��l2ݽlg��J�7��^�����U۝�먔lX�&���_nj}�\�~w���f0�������kS�ue�����D�ex!$#YM���Of`�{q?�i�7%܈��"���ig��6�!��J�A�}��;��y�D���R�\'F8���H���XA6�~�Η��ΰ�S�MxNAoIƓ��4a:K9OKʉX���O�8��5����m����xR�p�yʭ �ץ<�Ҥ��:0��F*`F���UZU�ś���r����XR0�&��m�$W�
3���k��j2{p{��2gӉ�`�)��'��U�3b,��}���<����f�5�l�����f��r�.^����tVw�%�y��ݖ��j�ע���C��uH���a9��p���`�����"I����P3u`�K�hY��Ȼ �yYZ�D*�A�R���I�W�h�0*��4-�<W>�Rp����Ĉ�xX��`��V�%Fs�6X���+m�d*�i��?og����-������/77ӫ����
���<[V��+O}u�*7�Z̮���j{�5Pÿ_W��Mf�v>��x�¦rs�.\1���l%�;7q�b��C2���߽��hW�F�Y���/�-��x��gt�GP��������#M��C{��'®~vw|[�%�8����%@z!K�4ˍ���RΈ�o~��*'l�;]_���ru��vG�H�j9^\�4-���Hl��:)�����BHޠ��$+�%�+07,L!k@������"C��4�%����'	��4�4mԈ� F�5����)��g!)�Z{�f�))%8����7sN*%T�Hi�DC��PY�$/a�s�	��9���~%�)ڛ�!�^��xBN��5Y=���T �l$ Z��kg~��B�SRqe��QC�M_5䜌��6k2�:-)�׈ǆWC`>��	 d�TCo�Ys��vd��ێ�ɴbr-3+Ȉ��)*&ՈB@C�8��<�z��*��K�����;*rIx�˨o�-�q[/��|($i̜��}C=��c߄�[�& ���� hN%�+ŢCJG�j�e3mZ��qY�R�1���Ã%JhNDb-X)��7W���&�XΊ����Qyʵ� 4VV���4Ɛ�6+�dQc۩��P��T�
���/fքrI�[�Q� ӑ� t���E�XƋ�	Q�LS�p��WS-S
��9�� �sZ綔! ��w��4�{y����g��x]���hy7O��\N�C�k�"��&�c(?Ǫ��f)<KEB�'��yRZ�'�p�s��Z!�w����XD�V�h,���x�Peǃ�CeF�U%�H�l�ݶ�q��4���O� �g�n�Hk���(��"��D� Κ�(�~�??��z=ΫY>�.�٤�EGH��&i5^|�lsi3�Εf<���$6���x�j���������f�H���j����_m��
sH�����,N����y���y� k��0�${�8�[�m��e�sZ�V���_���qÔ���:9��j����~v�N�w�@FB�D���pCY�@0'���]�52^Q��|��ڤ��H�3<Q�LS�!� %n;���72O���f����������wn�0����t�IuUB�N-!Vr�7@J�I�!��RRK�eTS9��T��t3�w��M�)�7E}Ee����sD�U���
|pn�՗QTT��RԷ�O0������ʹ�UW���w���Sٗ�����O��	�#C9UDsc8����r�>��pU1f�E��������*�K�S�_��&�gP�b9q�T����k��>[Ĥd�H+�2C*�H�3L��Rs�/�����^������է�/�������l�ep�a�J͈�C)Ԉ�-�DJ�E��J����nR\�����6����XAQو*a	5�[A��Y:RFi����P#.���Wz_�����k��o��7}�\����f���(��	�V��f��|�����^��Q��GF���`~�P��ܡ�=q��'�VψK%|��q���,87#�\�s���<)�c�9�Ŵ?�~� f;O�;W|�y��m��Ͽ�ݧ_��)��_|!8 ��o������@�M���XU�O���pgԬ��ӻ����I7���l����ח������M��7����z���w�a��Γ|�7�eS#�`?c�\e�j[w���|��wCU��՗J��{�_o_� �1��@�;��~�=�����e�䂱�TT�R�U�}����� ��Y�e��7ն|�xn��e;��0�g�^�'��m���RgYʲ0p��s�=D��"�G�H{���.�U��o1pTR�C���TX��z�})����{H����[�K.CEY+��?�Ez.��N*{.����1��#�X��#k�2J��Z�	h����r�N� �:��٠���I��[�8a����V桁u�P'ƳQ=���ŲQ���W�Gn�i������P�[�O֊�d���Qm_��r�V�l��2@N���P�x8����-����l�B�I a��3I��v��ⲝj�H��}|}@�ys_�SE�4q��x��x��-f��0����>Ӂ�/��T�&���H2���(���Y�UM�:i���C)Z�^dq��>d{Hw�X)U���cc�T;�)5#-E�~�{KEZFܥ���k��àN9��,`{H��J�c��cȄ찟�Yp���(֬8��-�5���夒��R��P��#�vdP�#lE/�#��#[�����ֳဪ#Ҭ���M՞��p�{P!�,#�,����CY���l�P���>1�<����n�k؏3qTG��'���,u\#�pO2q_��~��C��iW��Z�h��u�P�Q���,Ɵ\��$��9�O�S5G�i�A�d`��4��c��Q�Q`�w���(/V��a�e��:�k�*{*�qH�9��h}��*�qD�l�b���=���ȸFo�=��k���w<�ڧ��8xʊ��̣-�7ZP�@~��Gn/[�B"�8�mu��f�6�����!i�ٷe8������x2yS��﷎����ڣ��c�/W�N��t��������Gܿ��5�f������!����E����PK   `��XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   `��X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   `��X���a� �] /   images/43b8fa2f-aa16-4fa0-a6a4-ecf006c83c4c.png��wTS�?�FA� v�c ��Hh����*� �J��[E��(V��b���"j�FQ0� ���tAj�P��9_H��1�����C�`8�����3�Z{흇��wn?���_:o��(�@v�n�߄j�P�q{�������������/D��oS����K!����n�hO{������ek�n/�扌���@�B�����0�5ho3<=B��n����t@�a����9*������*����&Ooh����p�8���x\4t�R�`Y�p�B[_T�w�o���,x���M6E���r&�ÅA�XzлwI^g[,晁̈���n���_�k����ZɆ�&�i�J�)�aF^��
��w׽͐�j�-1SwS5fp!���,Sw�<�x�m�S?��mO��
�.|��Tc̑��Q�a�P?����-l2?:�����:	���s��� Z�E�����pu�|5����h@���}h��|�/9�Ø�'�<Řj���/O!ݙ\�{<$�A#��Ũ�!��@��H	�����դb��}���f�:?�q֩ez֬
�UD��'�.�<�-+Vg"�w�v�=<d���Q/6r��<�z[x�zE�]s�=Z�.6e�7�G�#�K��R�1;{�芜��J��њ���SU�@���8�>��R)��]����ak�)_�C��8H��-�k��yBE�^[�T�t<��L.S_JUlWU��`~�����K�.D��h;��+�n�a��Zk�J��Q��͛�ݲ]K|Y���`N��f�6����0<6�vC�c�\�M*T���m|cu�0A���9�$��D�Myׂ,�"Q��R76!��C�x<91�>5w�ƛ��T�SlR���+�f�5�ã��Qw$�j�]����:�0X��f��\���i�s��s�l�7�+9)C5��^��T~������<�:���E�"������Z����Rsؚ��W��ƒ�F��Y��f��ar��I�N�ٔy[&g�2�X�VZ�HH
e��zfDN,�q����3������9��>A�\�:�^m�K��W��r+�11)���nn��k'���"�`&*휶K/�ƑPI}m;&��M���U��i�gԸ.�메;(�Djg
B��	�:f���cT�HX��ѣf�\ʰ7?4���Jb1��_�c��w�M���R����+O�%V���L\9b�x�g�_������d���S�^_
�݁�d�vq�l*�PҌM�+�.�C�Zꈝ�F��9øcN�;"_��aS�K/g^�P�x�!��Aؐ�м�R�V�?y[�C��"��';�I_橏��:U,��F��^��� >�3��9\�y�����������^��2v!b%K;w�3���i�9r�ʂ�
_J<f�N���/�Wmi]��R�W6}�0�ͯ��#�5='�	5�c'��p�H+UP�Mֳr�
��DI�_"��ܩ��.h*Rc�D�&z"�~(�p��I*��N�>�讁�"�܌Ι yW^uV��7/=
c~ڕ�_��&����W�2�1��U1��(��n���j���� 9b���wX�^^�de���&�f��M�����W$4��k�����s&�r�J�ǊD�_��*Bvdb��,2�E�O���ݐ�+�Y�=Y��#��l"���}5�%�Q�=�ߏm��e�\Ω�B7�3�'�F_��gs\ɲv\YC,`�*3����hhg�}��z�y�2���v��_�}�6�L��!ˣ�g8�D��.�5�+l�s�#�D�q�_}r_��l�H(�T����F&�Mrҹ�&���H9��$q8�dlkZ���/�K�VOwG�@�O
S�C�΢�Lj��@�����;�7��034�t�A��7�8.į_:�O$��Q8� ��|_�e�I���5�Ώ�i���3�fʁ_f�)(�����m&���F��'���|Fw��9�m��v��PN�~ r�Ra��a�sVr�Y�B�7������L�D,+�kO�I�ƴvc<0��S��D���K��p,Ah�
�C;x���P�kcQ�O�a靲p��!���x���ѱ#�[�VM�/5�3��¼���!I9��:W���A�ȵ�RA���%	�����c�;�E�δz1������Lr�"� A9��\W���NR�U��=����}��/7�>?*���$�D�c�2��2'�cЁUۑZ�_I�p�r�5�^e��(��^~��yx��Y�Kx���2t�Ne��q�����O������kOyb���喘V:��3� �<�� ��kH���~��$���%~?qC�:B�i���M����hU/`��9Bm�9�
/H��;6V/U�QS'����<�6���FV|~<��1�L��ᕛ3�,D�
}~J��LMjF�d%k����-p240:ԾiWQx�Jc�8�G�H�m��ڝ���W?VW�#&1��'F�5Rnl0���4#]�\<���9?nI{s!�ߢ<<�Q�J���\p3��(l�\��Q��煋�"OxR�F�uB�����*�I�"���7�&��AlQ�H���p���j�����s����0V:���y�m���tA�I�s��*�ɔ?u�#��w�y�%kh�?e����=�C��O��f����0�g�`�����-p��i'��*"Q�`���F���%����JV.§��u���x��k�I���U� 6]E���ڼ��K��S����ȹ�B!v9Y$�n��{�G�Y�+V멷+7�|�C��O&�kb��ڲ��q���у7dI$�d:�+��?�ܜ��h���ŘYFj�I|8*��ӢK��8��3������x��z����)I�����}As%R�1�����z^����X�y���	ϣ�I��n �I��Y#<m��*�_��,�H$�e� �ӆ|�u�X��S�JVn�`�Y��CE#?38
J�^�<������ޞ>�D�U�a���:�IΧ���T��XK4��NI��ɍssδ�>�lY���S�-�*�������~��I���̜����/aS���d��#�5V���A�9���|}z3�k2���_�-�M�,�x��&΅���MkEۭ�n�k�#���N�wcϱ�|�\��>���JE�͎>ߗel\'����.E��ީ��/2�"IJ&�6��{���s�Df.�v�|��o7`#���TJ_̦�4��Q�mb@iO�W��dTf��O�j45&%�2����������K���]�!j��TWǌ���WM0�nx���D��M'�
V^x� {����;��!�*�S &WA�1��Y����`�C2Izf֋�M�z�ą��V ��,n�?�2ޭʘZD����mt,!��ꤸ�B�V���a;��
it�*���=��(�@:k�Q��M)�!=����@�(�r�{1$�2��i�_���LNr�1%M
��`|�j���R�3�b!h��j7��^h�^v��d�[Kd��m�Ћʽ�,�R(k� ������4b[M��wJP[u��k�uV���N��+�I�l��[�!/�T�Ҍ�I9��C?�h�<i��f�$9?�&䈪��aϋ:A%��֪	]�<��+���%&�WAT���i�+G��$"����Ȃ2���V�����z31Pf;��hbC��$�DP���y.!6?	�g� ���J�+�+��6~�w8Pۨ�,mû��8c���W��Z7�:�$��ӇZ�x��\p�~Fj���ڒ��ψY��?��cEs�X�l�2Y�膵c7|k��;���2�K������.��'5�9v�xe�.�4�]˵�1�a�@9-�OW�+�w.Ǧ����SS�4��1C!�kr��$��PQnTOtk���j0"�ȸ���52���,��I�c�Ý��D�#�1�]b�ck��/Q�D�
�_q�s�|���Y`�a��6�bl��v�jP���v"�e$���a�>���7�31�߸��eW܀���n�#��
�a�_y��D0��&�d���b��Q�'���1��d�F��Y�@��e&���aϖô���2�։��z�55�$P)X�{�u����4�aY��n��	�|���	�b���&Y����F�Q]�$�U��cH�߱��>W�W9�u��qn��PMy��LۿN�OCj�&�SW�t�/����EB%�]-ƀ��ߧ#[y�J>�;T)��D&;xqL�����+�"_�w��Q'G�_]�#>�WA(�]<���m�I�u#Q	��oECֽ��<&�i�8�Bв��փ3�Ա��KE���B/������JJz�s�`k�Aϰ��s�>�)Q���h^��1�
�+�E��ɬG�K��=u�_ΊI�8Ҷ��p���v�^�o;�3<�á���uTN�s�k�ql��]�~��<��߼k���y2}^p���W�*�O��`7"*��ޗuun��Z2�N���W(��H��Y�t�Y�9�}#���������@��r���D|�@u9_f�l��b�H�U��n�E-]C8a�?��*�`�q�t׆GeG�+J�aė�1LS^��,E���ji��	�vL��G��F�e!�v��0� ��y�l��5S��0�9#+���b�B��
��@mL,��v�C���yu�Y]�G��I���O��/ƕ��,��h{Gu�=��L��H�cAK�t�Ѫ4v�2���N��f��@7�@�"�A B���g����]f�����(~��^�n7d�"�A.=	\O����,}I�rŨ�ဈ�J+UT
2��R��#7���z��wn�A]��Ly�09� G?K�`�>�z�,�"�L���A���@p ��83+����|�P1'���~p�+�s�	�(9����큒��+���Ѧ���~j�Z�G��x 6�$X����t����k7h[Mg��::S_���6gA�7�j�� ��CB�������n6��[{�#�f&D�sSFcz��x�WؽH�3��X������V5�v�(�Û��IӚάˎ=_��eI=@Og���>\:���H�3�S��c�����)���S�����=iF�o��<w ԐZ^E�շ�r?�)A'�3/��rN�4�m��N�ж�oNI�߃ M儊�(#7��o⎬Yc����BRu�=k�%��uR$���W+�-6t<΁\���2)���s�n��Q�@�-x��h8Gm>�.fٙ-����z���#T�}�k�3o&�1�k���h��������dK'�%�e��ZF��-�c�ƺ�-��З���dg�kyw�53���7 �e�֋9�y�$��ˎ-��ɬ�@m��W��p�7O!���i�W9��xmv˥Jm�=���P�����8s/{�����q�$��x��1�qxT 6m+�sT��Fk�%#��N�l
v K��Ki$�-L@f/pC�:��ƒCQ���b�Q�}nN�Mj�R���C��\��i��ZR�L�el�/�>'ͨ�z�4���΁��!�r�_��n�_AG�Q$��%�Pu߅����L��Xԣ�O{.���cs�&�� 7s�1(��i	`v�Kr^g�E��/�ܑu
�C�����X��N�x�P����W+1�o���E�}�0��?����:�W0�llɪ��so��9󈅭x2�\��'.TUu�#�B?�Vk	�'�b�ō�G�--Q���ǣ�rP<�`�xLk�1��r�(�K�q3���&��7��]�d��kVWM) [���
�ā��Ux�ī�wc�Cp�#HT�G�5�1⁓z�X��(��y���f$�µ���Lz�#~��QMM�>�7����ķ.a�A��T?�53��5'�6d��s�.ܢ��T�F��i;�G"��
:I����t�ؐ}�� Dd�V�P%v��F����R��w�i��ENu/-Aך`wW�~�V?LOC�@f'��VWJ�c�Pص�=By�G��sG�������e�P���0oB/l��Q�]��;P|���yᐃ_R�LҮ2����ծ�X˕Is�n@�M�e'I��ͷ�AlUw��Q��d��"d+��O	`��K�n�R�c?B<R�e]-6Ig�<\�b$w����>�ҵ~��f=V|5fs�G|�-V��љ�0 _���-aCU�2c�Xp$��+W ��6&9�+uz��"H�\8m�z��mT���ֱ �`��{�H�L#���w(�/g|
�)&��k�E��Hhp+l�-;�)M���Wz�&��0�N��I��}��,��"�i�p�u1��D�D3Cn$��8�B>}�쾿��t�W�]�O�<�ߖ��n[�݉ߋU���\s����m�AQ`�o�);��_/�Kc��Jlܬ}����}Jsug.���]��ų�,��
� L���J��te{���0�Q�f��)��E`߻�̬w�U��]�2Au�o4 ��q��:�@���3��<d�U#2�.PJC�|�~�2��L���G���p�m}��'�R�G~��Ű�>SC����<C�"l{��\�H���>�g����C�z��%^"
�t.}��M�����������7(��ɱ��)�sHX2W�٬�����RZ�17^�������Ёi$��ޞ���
b����n�s٤��|�B`-�5$:r�V1P�m)�����9����&����9km��c��{���x����&�=�#}t�?\��<~�YI�^��q,�Wy�V£A�X��a!b�
?�MɦA�7ம���Ee֢��%��'��d�7ېYv+��,���F���Aڱ6�Zo�V4��>zƤx��k������U����[�X@��K��{��F�f��.��HU������2��˒�w06��t"�X���%+*��y��!�Ș\ۺXX��Ɋ$w��<䰖��@��������yG�Z�Cb���2r�Q<�Y�ʑ�/]�
�2�~=��2�fơ�sm*���&���6X�g�~���SN���k�v�!F}}�M���
�S�<�\�?M�,�:R@n����5�n�|H:��Tq�[�hj���s�I����L�Ɨ5�`��C�L�d֊��e�Q&��G������2��1xE���#�#��\�t-j�PW�b|8�@�t*=wE��'�p��63�l>���8��D�>*���<�o-Z/�ݸ�$b��DH@��{'�0�,A�E��H�� ����58$�P�F>���:$Ћ���C*�����\%j�Qg^�u�j���X�1��� ě��Y���.�ڸ����C���N�����$m�P� �x���јFv�{�Vo���2�~*Xg���P�ѓC�͛�Y��v+0`�׳�E��[['� ���-�7�&��0e}�(�� ��c���� �����b� ��d�T���T	4�e�8畋;��A���U���f��=�~�[�gF^=���|إH�F3u}!��� H��).Bm�QEl�x�%4��Qsx����Ee1 ��`��T�g���N�p�������x�7aP��[&����X1z~��n\�)�־yX���Ӯ_�T�0�/}<l�DPȷk9�@�"��c��8u?���b���u��G�J6�n��a��\%�Y�3�q𼤟Yy��Ķ����|�uUڍ�+$[����Y�{���lC�ъ���`%�Y�᳏ ޓ%e�T�+�F���}���Ό�G@b}��-�L�����
�ؖ���g ��N������5���y��� �=�#���.��*�&��7����=3m�8�`8�1����m���m���YF�~��q�@P�$�����s;��'�����nX�b�ג�K���w `�pX@�<s#	�5�f��/fW����v��klǳ�ѓ�U!y��>_/J����z=��_Q����[MA���22��A���r|����j��~J�nS�����'���q���ì��D\?���%�QAgi$��P\K
���+�A����r,�`�S�V�HVy���~]ay-�.�ҝ�����!ͣ��*�w�6&�ʹOUj6*���\a��zY�\�-~L8Y��P��e�ߋ��l�h����-�G�������O>Wsv�z��my;y��T[��	>j@#�����k�|����xLh��rb�.���$T�Hj?Wت�v4�쐼^�t��<xE^Zi-d��Rp��#��r-�?����N1���� 0���0I�w֛���0tǳ�h"�(�qB��c�>m���x|w�1`�BU�j%�ڴ��i��R�@"���!�m�l������u�i�A����kӸ��I~{6[\�����2k\Qѷ̓�mG`\��'��������x�@���^W5�p�2���_��}?�./�r1��o�����	��8�`)� �1�5{��lJ;����>W�T��b��"Z�$V�]J�j�ҋ���f}��&�VŠ�&���)g��x'�Z'��O���c�~c��Co��������/`�ϼވi�u���+Y�$b��ȘO�:��~A+۸(x4~��sr���7D�۷�;�?)��
�m�ᨶ��p�F�{�Lw~���a)@7��:~˩}W�v�W������G�N'l���}1�8������F�����5L���xw~"�|��ʋ��nl�7Ky��?����j�����zl�3�#c��ɮ��uk[!���J�]�o*RM���8[Y�9W��qu}�]�~~o���,�&j����s%_�i�!w� qmV��]����9F��;Z��r�X�(}�搻��66a�"��h����f��M��!uw��K��Y��Yj����I+� <Z���>��Ũ8��X���#��-L�sd� ����s榭�;�x�?����L0si	?�?���t�<���]It飔M^��EQ0�M���浾�c���W����Hħ�������Q���S�Q�x��t��|�m�?J�8�!�椠���
��u�R��w|�0l�f�Ѭ�Bm ~�m����$ȹ:�v2H^~;[�Hm��;��V�^.�H;P�葏c����s�w\=��A������\ �jo��;�, ]�A��2��d���8-�CBE\=y����ְ"�Yg�YH6��
�5�3�S�j@�}<$R��}�O�w�q{����R�~�w4@�q��;#&�/���(*��Y�v`�=�v�Tԟ,��ڈ#�z�݋ �i�Cf�4�?a�iP�vZw�c�	 �#����T=����zh
j��tݛ�������"�B�UEwޒJ.ǚi���8鮌���L������r�rj�ӭM�
��2����?��m����n�V~WYE4���֪�UD�a}�Kn ��u�r�:�����k/��S�I��b3}o�윲s��� ��y��o�����Y;P<t��3.�+�����?SXZ ��|�؍����rc=����|E֩�=�x ���t>���;��&���NN/ҭ�:��:2v>eʽ��j�^�dw;T%���T;�5֚#�:ch�]�0�1e�u�H��N��bB@�!��4�b�<�8&_ ����h� �um���.VCy�05��N�:�=ML��4k�m~~3��I(�=�� Hj�8�{e/�%`e�6/S��~�2�LC�Ϥ)�r!��5}�0i���A��ea���m���%�Aa�0���#r��7��r)���;�v�k6��&� �7�ԍ��!drA�k�p���b�)e(�x#=��jC��2v;vZ��{=,H�:K�Qv(�Fb�-��^ئ�
X�+�૵X�v'X��T��G�!
����q&�T�j�c*�X�5���#!rqZ���&���b�8�wP�gY��K�JS48�`����[��Z�a .�BH���K3������!������|J5�i�Gֲ8��C�	��V�M�6��Ok�2N�2�Y��+xZ��MZ�zb�W�X��\���tf��av�A��^0�'�����k��Bꜿ��{��.�2��%�ev��-z�|�so�Xм A�������𰳌|Ai����%f���������-���Ogr���K�
N���0V�9fVB�o2�]��.R�d�?P!џM��A8u�:s� �	>/�SNv��Ћ��}m�8��C���ZN�г����N.YÜTv�	_����]��$�A`�i������m��l��ެ \Fk���6R�@�kןב�����9g����>���?���հ���cA>��^�������Y��7PR� ?(��ͪ�8���DlQ+�ğfO��
���^�-e'~����㌼p�?���zJ�I�z�ZdW��]��������yQ��Ϡ�&t��Fg���1�@���2��8�R��P�T��9S��_���5+�����f38Ʊa��jO�~�6,0�M����5,*4�l���?<)94���X�� ���{}S���$2��=��O���rm�T�L���+o��=H(�
ք�����j'�	Dݨ�0��4��p�5�Q[��c����%���%C�!�5���XRن�E�w�S��3���<��]FÔ��{�-M;4����&�4<�� ""ذJ��C ��2����}a�J�$;�bz���a<X���x���%�t=�L�;S�-���~������G�8�7yw�쌷+@�Lq2�;��h,2��o���v�T�s�\�7y��L߆��*U�GM3��Q/
���MN�3��7A-�}y�s�Iz@�$Wmd۸2X�����@G� e�E���^��1T�=�������˅���M�<�c��~�e$a�@^����8b�ж~��(1�M�{����)���y��`�u�h�c�ʹK�}�l*P�M1u�7����kS�D X�)^�2��=.خ�|�q�P(	�cg��$ϫliR/��j«@)�))��*��a���N���Of8:�cϘ�.����9�񋺓e�=g��,k�c0Ǹ/�X7��b���� mIl��̍f!�rm��w�x���嫬���m/��o��+c �3��$?Ff4O��`^)�n_/L'u���3o�{�SP[��b5X)��l��+�kߞȢי= �d��{l���'ӇF�z}]h����~N���f����1�X7������2%	�'΅i(��������p��dW�3��RwV}�DP��%�t���e��2f�@'�)�n�q�<�x\*ץ�œ�j��x�s�T �}?��pk& r���bi� �>��p���4��f黝O�<}h|%D�]�wg�RX;���q���j�u�M�����s�h1���Rdtz�t�A׎�8`<����'��V��@?E�.��P�+�%�S$��BU��OHN��Vz���Ϣ�c1�@���}WO��X������Q:��.�?5�f}Վ3D~�8�UBۙ���q�3m'��L~[x�O�/9�b�O�ZәC����J⼙�-�3n�"�B�`I2�y$�>2-54�P9;�뾼����Q��hG�C)M|Ci�m�MjL�/e�ܿ*����ĄϪ��q�ng�K�ns��ä_���ő�s��!	L}!�E0����<l�ʞ&D�ۥ�R6�y�tX 2EA��t�h���$0K!����|������37��{�,f{)g�F
���AeڿD"�%h}�A>D|{U^���	�[�����������Hh��Ao��
*��#�&[b˨f����Y=�v#������ʠ��C�jX&ca���
���DX��ȣ���^.�Ù.��-�G��
�!c��q�s��c�*g�����y�k Ү�=(�`,�r[�U���j��%���z*�]����8��9��{�K���+
a&�Lj���ڭЋ�ucg�Ԡ*��=��������
	�m�G����FA��n�/��>�Z s��?4=Ͼ�E�P�i��>+�V��-0�ԯ�=ivQ��`5|��]Uݱ�NXE2�[D�!\�]�l66��|t݌���.�"6���g#lH�<�Q�ڪ��x�E1���m����b��F G; ���]\��0��Ɨ�z�Q�1��V��!�~X��/k�>; �-�G�����4Su���F���!�������
��e[��j�L�,��,�h:�b�)݆�$_l�j������Ӊ�-kw��UޠS�Y��B5jb�Iڹ�w�h� �KM�2��x0?m���2I��}�-<�j�x��e̔3��p����C�	p8�|�(Q�
��
�O����-�P��Ue��V,%ziƂ��/.]TF�B�#B��{��&��60���eG���e�3����Y=ڑ�v^�y�p�ߓ��Ԙ�Ս�կ���A9�Y�v��"'5�E�^�S�k[�M��Ӽ���ti/_�u)mPW2�.蛅�_ m*(xRiv��}�{��n�?h�t��խ�.l������+�򀂂&#ts,�i�%�������<f1A��l󑭑�-fǙ�Fu���g�d7���B�!5zW��	 �z�H�g�)��:�$=c2�be�7Oi#��~���v�R9�fB��kxEj{K����]��m�hP�ˉ�K�fl��7��E-�kRa���.j�]��6c2ï;�����q�l�l4�$xb'��<�(�ޕ&B^x��s�$\��>V�Eg�&����3��I#�^��ȼ4.���&����Ӻ�Γ�Im�q/�lY?�Y�p�|C�|V�O/:�{8�qK�N���yS��O���t5�J�h�vߺI�0I�Y;8�����ݐ�W,�l9�"�(�_����9Ί�gV��i�v0)ǲ� 5[����U`�6ȃ.��I�Z<)�k_���L���c�!�75�����~g�Eű�Ú�T�����f"�-@_���y�g��ve�`=��a�$��3
��os����I��ys�`ܟU�D�z����L`�__01��7��y��g{֩x��s<똕TwL��Ϸеc���.�C��0)��3\���zsJ�F��*��>�]��I��q�c!��'h����Hufiāo�K�yz�@ ���=|&�� mH�����Ig��c�.�WCDM_j1�C5�;zi���z��x~%��-�imK_mN^5=rr��B��EӃ����$P��d',��1�$)�"��`Q����d�}�委c}�H��P�s��_V�S��(��{��s1[H��!�ْ�ǅ^z+>?yc>_����L��#6;�]D�)���i�.?��M�=�,\	U��˩@mW�Lٳod����9M9�����TX��eCY����6�g]E�Y�9�]�nbi���+���?�ދ��.���_�	�F.�[�����a<�㙒���Ⱦ^�lx*�ZG��&�V���W� �hdd��͂��<2�I�$'�C��P̈́xF��.ˎ�R�/�� Ƽ�%��5���>�.Fm�*�X�n@`f����IR��1�j����	���o��nO���w�s����#�p�����d��]��vz�L<���%�>a�7&�_I����d=��Z%��0� �<A]�H2Z���TA9��i�g��_ f�c�)I���z�с̃�n��I��3X�p�A�C?��͢��bl�PWc���4���"i��L-T���TH���cʓL��\+(�u���:�$@�{��PՖ�stj}������v��'�JI7O;�;0^��z�	�+P[��E2�~��`�`E%�G�]�]����7�lLG�	�,<�e�6�U+g�n
�&����|]<֥�*�������Su 169�����`4.k�3.��o������]7ӟ^8p���PU�&I	G�(m�g��N��M�[g(о.���{ؠ��x���N��7UDM�j]}_��g���d�E��eו�:ι�4;�o	k}�jI�q-�����U]~`D���D��5G��,�u8�vC'����~t&��/OY���I�5=�5p\��2�(X�'x���~��O);rw �U5�nx*S�ӗm���a�f��:Tg�[6��κn�&Uz57��i���t���.'�t�ԚZx�iqNu��l���'u��+u0 ��	0�G����.�H5#��������p30�(�RN*����9h��E�Lr�ڗX&�;�P�F0�9MK+5�1��A*�S��߶��c��.d�K�_K���vdt���~P�F@_0y���v���
���X;L>�c��&%��q�ʄ�	�M��U�<�a�0G�a�K�D��2U쌕�L(u�!t�l��S-F�����Jg3�j3���3�	7�&�h�l����aN�r���{X��$�\&����!bˈF�~��rb��y����у�'�3Q�Z��}��N5�c���M>�ˬ�@�H�ǩ#嫬կE�H�<��^F��?
� 8<[�
�\S�m�w�e��,� �O�@%w���j8⹵l���h��;���H�ZL�$s͌w�.6қ?���cg$'�r<*�2�&G�+��,,�'wֻޱ1Z�c�)�W值�V���o�VS�5�饅��HV�5G}"�0��б��CѤ7�Y�c䪗�<��V]˯tn�CT7�ޘ?7�5��������Ty1�A:+����	7P�W�PW�-Kd�L���@2E@��(I���!9��<ITl�ӝsv�7h���7�8G}w�~��2|!}��d��vZ4��<��Sk�)A
�9�$�Ѯ���h'#�rEו�=��l�D�I�-��XX��&�9{G!e��7>�t��[�5_6�uD^E5��LmH��_/4�Z�U��5����"1��F�:�ܣ��Ě�#,s4s�$Ӡ���w�vE%�v٨e��t����3�Ip������-�Q���wB�{�'�K ��_�$F��b�
d�5"T��;u�����b��L�P��5z_0��T��DEOa���}Q%E���V�Rkα���pR*Tb������0�5
�>�,>����d\8}H��O%?�/UT�`8��F@�E]$.%g^�)�nK����=]pxb�`�aSy���X��O_t����<*S�ҥ%p����w�e��|��DLܼ䍤�/V7�NA^X����1�9����eL�~��l��#	傩Y������n������������Ҫ���0QX�Q�7t{�Ji���h%��"=q��9��HWZ�����\�K	�����M�}� �/�0�����__R�����S��<u5�g��������c��5MC���~Ft�u��� N������Z�-�� '�Kr���xf����_^���N��r�2d�4{�8�����7��3���7��3���7��3���7��3�?�aU����Y���3���_�' ��UA�������\�M��i����3��m9#�6w5���~xk:�{���mZ�����_�:���Tj���G+i̊����4~(A���m{������'xי���c�m�N�ף���ϴ|BM�q���J�{N���x����B��sts�G���v�9��V�X����t|�dPEie������ ٕ�6�Ʃ.��/R���T���_6�v��϶͜�Q��3�o���_^���o����f���o����f��Z�����-�����\KGB����g��>�*B �Z�s�=Y;�0s�\�n]"d~�Z�LM�!
���sp���B���9yv��%� ������n�L�.�3a��A��f�xJeo�)�0�Fb俉x���ڹe���VE���ܣ�ȯ��H������|�+�|ۨ���3ǧ{�ƿ{�M����4�B��P B�]��~`�����^xy��:ǯ������O�L��j�#9�M��7��sAqS.�}~�ￇU��o�II�p�����G�����\�s��7h=|(�4�/��l?� b�5��x�_��	��"�T3�Vn��bw����Iͽf�����z!��O��N�/\t��x�O1Z��r��=�V ��r"Y��R`���9�H<���Q@�.+Mf�����,[��-� ?CNq�m�[�{�y~��2����L���п:���6�?D�R0&g���w{ (H�&�E��J��e�H��j��Z��Q���#��)&ƿ�sS��SSqK��-1@dw:��G)N[��rRW�3�Vj����ã>ICl~�)"����3��aF���|�Js��`�]�(ч/�	����x��uY4����z��n�+5˥��ݤ�-�I?a8���V�C1��[��)�����z至=ʻ���O+�Y�L���zB��Ӓ�Ik����?RۯkWE�<_Y�B)=\=�$<�n������w��*8�;ikf�2���'D� ҭ�����ә�r@;����+u��ϡ���q��?4`�헭?v0�`�y9T?*ν�j{^vP�M۽G�[����Pm	�V�����J��]���;�Ŷ�����?W�6��[l�g��	3�HZ.�qj�> _�q&����5�E� �+"m�W���i�U��7�-S+�5�NN�>5�x�!
�~l	�v��NTQ�xD�
?��A�Ҿd���:r�� �9�ag���-χQ��7�|�د%��� 9�N�!�m��y��E�_L���F��H�)�뮖v�*����z���-�t�����峇�>�<���������:�GJOuo�UpO9���j�<���[�w�5�)�_ >���u�̈��5�eK�+{敮]��~����ի2i�wo_w����	�}1��jr���~z���399�������X�PQ�c��c��QD�t����?�� �����F>߭�ٲZ�=t�|46�G���e{��9t~�4�T�^}��e�x�b���6�����h���%r.�G�ɸ��>�����y-h�s�b<��4�Ҫ���k���~�=cg������l��[V��ͣ�z�P׮]1�&��L:j53�g|�О=Ǝo_�%C��#���Ll��ONH�z�W\�oo5&�r�~��/;ʲ��{��X�T�8�x���}Zݩhl����=����-������7�mds*~`��y���T�����W���:``����@�T��ᤊ�z K��K]EAC_���umñ=����U�Q��G��z0���%�T��Z�	�O�3���t���ҧ0�2��0�@�	�z��6�6�2����g�]t�բ�������G w��&�P�����e7}��2Ґ�i�s�Y7��+eG�Y�>k�m��i�=\�J%������35��\pke�z�t���?Bs��T}�����t_����|ze-]��);�?I�2z�f^���Dk���^�[L�ٶ�$�s��F�A�Լ��RRF����CU�D�=�W��~�m��su�G_���R7�5��*��-�R-��\�s&��?�
�,;�����G�̥{���%2��f �Ϗ򳚆^���nt�f��Z�#Oލ?�)������?��/k]��K�*;�V���+�N,?�%��-�`�{<R}�jC��/�������D��2P��KA@Z��K��KT$�< � �}��C� uh���u������1w�������3�9���޶�W٨�՝�ت�go#�th4��<�l��^ Y����o�n��.���O7|�;r���)ILҳ�p"_"�ɉ"9���;Ƿ����`�o�ن�����������M��m��i�üʗ^��ϛ�b?y~�ӯ�Aڕ�x|y�S_��L	uY�R��{��mwx;��-8�Ms��dPaӆ�άع���\���up�.ʜ':�#r��E�.�(�b3 ���?�D�m�d�w�<�hIz�V��V� q{�t5�����4���򞦏�.�W��|2��qa��� \�+#=��	7ab� ���	�k�"z��쯻G��h}�Vg?���&y�����`�}���J�Ҿ��ł��,�Pj]�M�0��߄��ܥm����!X��Gi�g54�ק^'�s���aAF�w�eã���𪎕:�˨�Ʒ�di�'�+��ֻH{�ps���|�|r\{��4�$>��
�tn�]�{�Xv��2Ť�G�c�Ey�Rh�I:�ځȃ�0R�"����u>%ې+ԙ*J'�ތj~��/+r�vH�a �pϒy��bu�Z�ݷgD���K/37���/p����7a�m�8s��}�Y�٘1���1���J��'6��z�>�H����",��H��#u$55�?���������El�J[�T���+"�O� T���x�=p�'���*������gmz��+V��A�a��$ۙ��.	^�U��7pM�����ĺ�_�b�0B[^�w��㯷])Zt����ik�;S��]>]t�-'��eZw�Q��|L[�6�P�v�­�@�'~N޾;�JGw����]��yOo�?I¿�������'#�I�]� �	Bq��d�G2T"}��miN)���N���$\�V*�zp�'���W��^�����7�D[/�΢wq����耇�L�.V4h
�S��S���>R�A"�E�~�5��ψ��l���	��%�a,�b�]�����`1��@�ˊ����\?jbJ����裠?�Ȓ��j#�V��O�2io���y<a~i�U��rv&�
MO��*��+�v���u���*!�]��+��֘u~�IgŖ 'u+;=w���o���8~{E��>��-�O͖H[����2 �{��+��L��n�Ǻ��U-TU�w.�w;j��8��þ��0�ĭ������#��v��	5����$�J~�f�b��7�-Ҏ��������4���54&vhI3����cԫ��_�0����K�,xbk*G��O�^��S*�Z��t�.ۜ�_Q��Ý��?��o��j����g?Gm.D�_�<?��$�~����j�s��E���0��.-�ɩ'�̌y��2�D�
��U4k��.��aG��ZFQ�����R������W��{Q�,`	Ro.#�s�2Rl��da�6^.ZU�7��В��" �)���MluL_���fK"��ew�d%W���-�툡Y,�a^���X�SV׺�glϟ�	�2�}��֝�����s�a���we�s�؝���y>`#�-���f��
�v���ޢ�xb���)�pa��2Rr����1��ĳ�x|YQY��ǃ�\�՞
�#���G��l��NF���2�p߂t�6���B$���wT-��Ԥ�����Ѵ�2r;���"?.���Ɍ�b��T�Ѭ���?�����庵��d�T��<��� D���37������ 	�t ��ψy��(����9��C��hu=�o�I�s�x\�}a@�� �6qe���������K���mm��)n,:��)��F3�(M���OG��r_7�`�p�q�I���$G"��$��h�K.Dʹ�{��:e$~)|��%M�[b4$��/_ֻ��?��ES�6,#@/G�$�{⿎g"���o:@�x�M�����{.%	$5��z�^M�g�m:�q�Nxa�,Lݑ)��O�0p�r���h�R0�vʊ��1�u3`{��������0ҩJ<i��O�A��|�se����l3�@���Q6��pW��D-�xA�@TOŃzg��F?μ�(����]����ּ��B��cn�-�eX�){%��2��s��lvV`>�(O��6�콑��T\H-#X�L�t�tê��,!,�,AqSVv���%��N:�~����r"���L��&!�
_-� ��t��p�n��0��Z�H���TU_��F���v��&�){+�߿����~M*��Ɲ�U�9������*��j��S	t��3Kf�4ޫP��88!�4���|�0ĝ=���Q[�,�3c5��ɓ+w՝1���ꭦr���>�_��(�:�.qe*ʈ��������)��"�M�d���e�^��4����.�M,�ϸF�>՗��ʡ����@乓3����)'S � ׿��{���XEf�
�f�yĢ�%�� �ג�Z�"����Y��&`pm2��>��:ܫ�6kV�a%;Oi�l�Q,�Z�S�7D>cbRt�.G�UA��s�=�R����)�(�ϧT���̪_���Yi��(+O�[̴�/;��z��t����l�5�R�-�����9��?�މ0>09����M�:f�6�V���i�"�K���Q�Z��|͐u����n���7y���b;�s5�
��gH��T��6�ځ��\���	��L���\J�t���W�Z��B�����;�(O��R4s̕*	a�M T�t ����ʛV|�$�:�4�x8�d�pbJR�M	�-v����͔�l��`�1�:\X�o��L�_�t/�a�����{�,��4."����:E�h@�t�"��G�`���<���3�+,Ԍ�Ey�_y���y	�4��ED]K�����/+����d&-顉��L����Ϭ9I�����"wW�Wɍ�pl�u
�bd��wf��D�QPbu��JMg#��]�7�|��ȭ�Ti�vW�R�%,]�T!�x��&� �O����f譁㚲�%���")rW�Wl����41ޏԶ��@�y8P`����8J�1��$��`_M�F�#��q$�ǝհQ�o�̀!hn�3��Q\pT4���_��8/C���]3_�!�IO/z��tg]o�"��FV��S��p3���jྋ�$��Mh�a��lb���ȵVs��'��w��ǯ������"��T�ӺJ֕����=��)9�}:�U�	��l"��l�tX�Amo>��|���M�;����%�a�q���V/���j(P�cQ�M��?�Pq�u;��q�#�\�`PK�'[�Q��欂;J����i����6_]Vy�QV��b����aHI����V��6�Ar�w�rYZ-Q �a,?IH�Rw��U�ݟJ9%!F�5�b8�#d쉶��u��F@��>8W�[�CSsIl�r�Λ^h������21qXx* F���F�	��a�o�ŝ����ϫ`'�:�[o���qi]�cpđӶ����M��H��fz�M��M��h�n	� VBΛu�<�^|���h�o����ޙqڣ�p�O�����e%����1#���8�.T�`B�0ȀH=�#v�h!�>ծ�4�i��������T���{�(�&@�f슧7v^����1�(�_�W�����p�����AD#dȱ< ���
E��EG5�H�����*�ןί�F��`���� ��7@E��Ti��F�-�+��B��?�v��J]1�G�SC�,�
E1K By�a�z��sܰ?�]Y�Y���*�}��������5C�ڠFk)g��#mZ��)�7_��Ѕn��Ei-�XԮ�9�3�j��p��a��om����L��o���:���j�W�ta�/�fy�*%�}V��:� ��H�I2�S���n�Y���R��bƏ9u1j�f�RI��j*(h2EKx�f(gDR;�T��j����QC ����(8�v߁�t�L���:�~�u���o&���y��i�xĸ^a�K��� 7$9П5�����iO�)�5�x�'N�����p8�]�¬o��P��(&�TY_��Jj��5�T^�5s��i	�`U�#��yӽ)���@�3:D��E�U�1�c��=��lm�D�KII���q�것k@pv�S��	�&�Ux5�(ل�d��KC������!���� �l��+�$��.u!O���ɇh��� î�e���Qֈ$��8�v�՛Cp��3��O���"�6Pb��%)�q��+�&ۤ�>g3��no-fϿ2���p.0�Ū�~��n������!�7��������B����Eۈ_+��ρբ"����3�!}��o7��{�y:�zq>$^�G�E�[�N�O/WO��=�׃}鮢�������k�5ti�Ǐ��W��N\�s���E�������/j:�u�G/����u�x%fZj�,��Y�|Y_�3��S����g+��o�4X�Zu�&�YA�h�=�H7Fv��&�Q8Rxn8ێ��O�ik�����l�Y�[h�?�p��)Fq��5^��JdI�} �^�⌴,?���em3��p��>O�|��0�T7��T8�Bc��`���K4�XMry�p��z�%1��#���9�cb悧h>��Jt}�F���?�ߍɤZ��^>��aR:,$EL�>��!�B�ɰ�A薦�nVa�V�B�W4z\l���-pzIn_9��x��I���?w�9�v�� �b�b>B�ʡ_�@��i,[Yv��Rs�I:��WZ|�'�F�0 ��M�OU�ޤ�U���f��U֖�|4eLBq�Z�#���VH4�]4���wB�ޮKN��U8�F�En*�	�:��婃P��7�11g��DCC���uPy�����K�Q�Pj�2��2p0��#I�����2	���,4)l�o�M{��+	\�G�C�3.n�[���k���ŕ��2~}�K��N+O;]\���L�"��3~�\P}t?��(U>�B6}�d���	�z�$��솛���뙾��/tYQk�̄�J-��۞�k>z��u��bi�Ⲯ��rv�#��3�%\��jpNT
~u5�9�_80<����鬺J�1��?����rݍ��7�6�I\eK�ʏ�3�ji��K�#����-�^��@ ��¡.s��*�2�����eu�\^��^��dDP��G�T���I�)/e���¬�3�Z�3����741�q�Q1�Q��K���U�6��@��j�\��Z�k�j�������K#�����h��B���p�~5,w`"g��Po$4�R�X�g� <g�ܜ�{-�y_FwX� 渘ICA�{tZ�T잞QT�n�X�%� ����FF���F�X��O�-���K�𐰚T>��B�3W�	7�p�jx�E�wu�����! @��}@���|��������/��|��{xU��3yn� �|4�Z1�&�}�+ /���h<�rչ�+1E�)@�d�Lzd����.����F��$$��[\�|�+W�y�H۟����*M6��U��k4�׌��4�Mbj�#�З��MCS���yk�e�5��%:�_ONL���&7f-��%�6�M����yH�!$���BSS=R6��rO�j�5v;o��ҝe��gB/���x��"X����rǀ��`J����u�ї�̝ww��:d�w{���˾�PqӯW,���h�}��?.�X���O��hO�7�����+�^�+�X#;�������e�2�7�C�1�$��3R*�!���*�K%+��9eDLq�pƳSgܴ�V���>��әP��	1v�:�Fq�v��.R|�x��AN�i�_%p8A������k�>x�.}� '�d^{%���㺋�ܘfu�l���(���{&�]��̋�v�*E?������70Z�	�ߑ8��V=*��LRw��΁t�<=����yz�y*a�� <Y�$�]�`[>�|Z8�i0���8�J]0�k��=�FVQ)A��f�y��(MQz&��:�.������aﴧ=�B�".�`b��B�;��r
���4��)̱������5۪8�N�D�3�5gD�+�ӂ�}Χk����&��b;q�n9<�	�-�����;N�^��,�-�-7@w��˖￳����'up�6���p}�˖��w�Rt�\����q�}�N,9]�۷��tu($;���J	SEQ���A���P�#8ܛ��&���ng��~����uE��>�Į�#�m11i}���^caz�Ǣ�i��5�nw��a�4e���,��NL��'"`G����I�nu�E^���������'݃_8y��ޠ��CS���f~�k��1}I�D.m��p峿�Pm5Z�|JdU^m��ZW���Txn�k���nD4,�@zW�ӏ��
�_D�/��/�"x6TPR{W'9����̯t��~X�v�(�y1E8�d.��ih��K�s�Uoo�31�,lnxZ�Fi�[�6����-���GY�{kz�������s&Hzwë�3����A�(��L�H�₂����_Uv��I�Z��B���s�/�{�r���3���A���+rb!7�����RO���A�ԺW&%��=+~����-X�wEVwP#2��&�C�j����ǳ�J����Geb�q��Yg\�/���"ϟej���Γdb�Ƌ���;��y��p-��e0�NrY��ڍ��έ߱�@���Hl��XD� �s"�J��%�,��|�����>��i��]66k5�	UtA�3�f 0�����fl����v��C��x�my|����Y��D�1q���8��!H��x&�7\�)�_X�~�5�-�KK�xӋ�X�
 ��2~��=�r[�&�WT>��q�ɍ��-B�[�?C�Z��&:;��a`�!`%ι*�鷮���c5O� ��ؖ������e�5��U��M_����B�q|_(ڿG�|tY�v�<�ץU�߱�	��@�i\s���B�0Ƌ��2�"p�S���.:��L��O�<�A��=Į�A+��k���>+�R��[*_(�4���N	�<�P��>�s���Xꀕ�Z]������9� #�x����H�7�|CdfT�{k�Sȳ.)��"�V��EM��7��8~�V�Y���M�.*��Q$3�m�lxQ�79�/ʆ��=��M�Ri��'�ӵZa^L/"@h�����;�_Ir�iYv�$�Ɍ%4�jo܂/����YF�X�(ȬjE:c�cQ����I�c����sʞ�+8ԓAV��A��X2�R�X֐�,\��O�g��"(T�x���G���k��@�>��h2��A���Yt��q1�����	���B(�8%�W}7��{���/nä��LG�k�gbo��RyԵ�;�� )�*��	R��q�5�}i���c�')�fU���g�������#��f\��RM��
�b��"��Jz���� u�4

���ڱ/�����\��@~�_���y��}�Hc�@"�f�a��z����M��/�P2/0'�>V�Adg��t֬9�	�g���}�;V�c��C��Z��Ӣ��+����x(�	���v�(|�N6=%&__��>�Td����mY;*s0O=�"y�paђ�蹞��% �vX�`P܉}�O�l)e�ο������$�y?��P)���k���$xO�@@�l��oa"ļ�Lͬ *lY[��sO�}�����~k�~���ϟRS� xg�}~� . ��
QN�Q��q�׺�I,�F	���n0,�U�S��^r��X�n��>#BHŤiG���ƽ�Ìo��>�G[�ʼ�������]�x�JF��ܯ���Q�!p'���8Yi٤`?>f��p���
�Sx��r���d��Q��;����3]PH^P�f�%)�����@���Z�TQ����0n&�x�G�c�p'�\���K�v7���.���╥����o�� ����I�.�
�vTo9�m���<Y_4�~;�F[?�����!�Z��k�uEv+���l�H���"���[5q�E�;�B	�CJ#V���T2��tH����](Ts�|	�ũ<���Q5盶�$RpFc��v����|�1��7�E�M��W\����?��~�~|����I��~���&;��������\���r>�:0�ܐ){A	�����B�i'�!%���m�J� �e[�K��z�M&F��JNSֹ��?�`�)*�k*'�5g`�w������+$q��l~.p�rc%��T �^!vAX*�x�M�LO �/T�����.%`�A��ߛ��hJ�8� 2�x.��`p��~ZW�'�p!p��F��pݾ���H�؅��8�I�h߯LvV ��EK�q�J�o�6�&��=�/��z`����a��W�63��
���Q���`�[�J{�ga��?Y���l��5>?��<�%H=�+T2�uG�ͺĘ$ �;�~�T\�ť럵4��ܒJ�.[����#h߶�^;���ũ��y^p�s ��3[4:���8����ԯ����77
���#ñ����ji>��g���JG��I��Is�4ޙ�����W�:\CXE���Z�����I6�R�w\)�jۣ�%�����n��j���G�z5�Ъq~n��{r�~`�T��_�z�3Lmr��3�|U�"��|�P��2eR��;�8��9����O�V�$d�2�˜����w�\·p��\�j/�Ių��P1t_�n���r�P0?���Dl�5��$�xx��y��"D��?y9%v/�^u��/�]�ng'��J��Z�V$y?9Iw/�W����?�L���j�k�5n�j��	'(��[�V�L���W8���}-J�JI����EZ�6! X�p��h�J���u����� ,m`��q��qN����4���i��I���[�&�U#T�\��]^���|���i�A�p��x����k��R�ִf�����Q�s�@Kג�y<��~�����ĘX���sa6�V��v�~OG���� K0�X��[��X�v>�# ��6qhS���Y�h���)�N���&�O���ZRp�tIj]7�X,L���Ղ����W�'�Q���덪���+*��RW5	�gX>�C&�<�<e�{&`�r�l�ڗ���p(mRğr�p�C��/,��egpM�ȸմP���u�/H�nI�`rҪi���3���1 d�E�`6����&h�>1��wۏ��<D+�/!4��rd�E>�L�sU�c� zX���u2y�!� �R\��4[��vV[��d�aMCd���Ɨ%O�9V���6����h�Z���) ���4޳�ʻg��t�t��$���4r\*CX�uݾ`�C�%@,5�M�3
2�O�? �K�LB��!*�eH���cc썐�9�J|�EN�Օ����l-vl���c�@�V�����K6�8tYd¢��iZdݏ�u$���W�d�)E�آ, �	Fq٦��-l�NB�k2-EOƪ�9�*��b�B�L����[|����De��	nI?��~��ޅ�_���nK���2o�҃�n\�wxoȇ��,��ؼ��{CE�*+�!,�s��|
�����S���C�e�UΦ�Y,�0�A�I�����%ƛ����5*i�Hl��7GE�x(J����._"S�ݰT!=������ڝL�0�X2)އ��G�Faץ�$�������~�ʎb���|�nᲈ� �e_��lD��n$ީ]���:�9�]�L$^G���l�6npȵ%��'>�M���m��C�d}�x�E������"PָX����h�Rg�Ӫ�r�G�^��� �s��'s�c�WלT��/ݸ���� i���T䱖ʕ���|�	���aϪ}��(�!�;�(I.���*��-����x��$���A�V�{��( ?@ED��0F��`�4����!{��e�(���>W�N3��A�<
�,��c�˟�`��@BF�Mo�,|�����R�+U��κ?tĲ��;����<�Y. �ާ�g�=�߉:yL^�|pF]�=� x��md$C���o߉�������_Q�cV�ƞ�:�$�1��8�P���"�|؍�-�Wy;Er��\����Ξ��T�ƹ����n��.�n��^��"@���0�n�*L�[�J{�Z�=C6�Z7�����+`QB�9U���|u>-ܺ�T@68����G�A�q{g����cE2��ԙ���~|�׆x_ +��C�ԍ/���zs��L�.'	ݳ7W�Xb�2^��A|6��3�͐̉q���$ ����n�ck4`��w�|����7�.��	����w�����2����Y�s���k��Kv�Ĩ�3����s߻�.�ۀ�bm�?�O��q�סHQ�	!@i�["�a��\���x�{�� ���!�T9�͜H�7�	_���Jn�eMԶ\ӑ?�Z��d�)����fXl�(��4:)d�6�f��Y�^�8�Z4zq���o���]���֌�	��8�\T����NI���c�"i'� O�	����8�r�]#��n!�������Q7��0�f�������.����"�Jl�_N���9Y�~��L
����bB���U<���k�<2���$�\���d������c��Dw�]�������R���(�<�s6�/�0�ݦ�H3䇊�3J2�Ǥs>?1�F�Ř0_�3��n_P,�UW�y��S��m�0�w�
Td#A�M�5��A[ύ�8#�=#��tF��.����!�WA��;:�ƘN�����#��[��V<e*~��K�Z��hު-���f��k�~�9������3��|f�E�~������cS�[!0Q�J���(�Ѥ�&�db_8*��]W8�Ì�����?�����w��I D�W��F�oّ�ap�{�}��G�f� �h'�ʻ�$�'`g���j�}�tPp�d��ݢt�����X���b�s*odQ�m�5�����*C�0Hro���k��D���/ ���RnS
�ӱ �h��S�Pq ��=�������ǥÙ�����%� ������EA~Ӎ-��2�+XO�.�޹	�|s�
�#p��#��D�P��mF��a����ͨNv�!.�T�;0�w0��_�'�|`�3���F���ɟ[���܉d�c|'R�ti5Shc�5P�<�3�����lk��h��Z��|���i����}޽@��4;a�W��4�ԏT�upa1h���f'�����웲���q:Ѥ�ܝ��Z��q�
Zs�p��aIԟ�IMN�y&Hu�~P��G-fϏ%w])����I�Av?k�{�ǐl�+ND@.�u��=ax��_?g�,*�k~�v�^�g�*�㍖߈�邧a���������ò���#�ψ�Ty���o���H�A��
6s���먲��~6�ԆWTO�d]Q
_��:��	K�����b!���:a;�ЎO��LNϴq	����O�SN�Hl����`#�^�]������M�$���
��9O�߹+KMP�)ꨢk�q�[��Y+#:cl�_cb����jg��K2�Z<��`r���q��s7���S*a�pl����'��^S��e�C(�3y�����8�ҰtOz���)F�s41���h��j$�fXT1�N�K�|�z'5w�'�H�drR����]�޵�k�b�X'�6 U���L��>1��G�vI+�lQ'�C%'t�*�w���w��P덐Ƣ\(Ti;CC�:�'�(�1?��f�W�A��<?ZO�D?̚U�\.���{T�X������J��Z\l�l���H��N<f���@�ٕ�Sɥ��P�M:�ȏ�p�����C5]<P�v�lv�C�|6��rr��΄R�FE�{����A� �����sD<���YR�TS��Y�O��m]m߫���K{hx/ >���D�,�u �x�[�j�I����$>���xF�y*^D������Q*��F�+BG?ͮv��/�#��Zh��;R�� �[;U5��l�}�xi��T!c��q�wO'(.�N�dCR>�*�G����)��2�c)G�ч$��:�l#�@����!gQn�Uꇮ���)�d�^���n��˰Q�U"ʫK�~|ʛp"oZUM7���;C$%s�5�#���bئ�Py��qm��B}9���%�35R58b'x&�"�_���ʏ?���gg��4���m�y.������p�T���i��>�/�BEc��M^ (�Ff�e�$�+��O��n�{�7����G�l�t�2���x��vɞj����EU�פ�X���n�c��"���f���u�tk� ��q���z��G���}������~�?袌n5�6�GJ�r�O��A=�DW�)ȹx2��`��e:ͽ��RV_t�����|�����4��ѕ7���/�TY��ږ/P%���H�s���3�N_�1����7�^�e��8Q]y?�io��l���L�[�Z�fUyaðqT���g��}���Oo���t|�[n/��)$c#1��K���kA^�࠼�o�~�[!ޥ.s�9\)��|�t�\�%�c �
VK�u�a��ʨ�� S�B���O�P���3LL'��Ԕ���������s\�:_Gb�W�S���j�����mR������-��p���.�-9�ώ��G,Hv@ޡ���M�u}�V� ��\I�������'�q�D��*�|	 Í��`©ca1���A!O���rˮlS��v���~I�*߈:>��OM���5�`�)��ӧ��}�Su6�J��U��'X�\q"�\�':�d�0>Jб�ù���t���PYqX �+_��E]7�(k<�Ll�N�l��cfHW�����?Xٱn�=�'f9yw�ݘYT��c�7h0
�@����}�W���'Α�y��V7ì|�gd/<���-�Qr!I�UY{�.�0�n$�}?cl�Y�V��tϗP�$����X���OϦgZ�X���1]g��ۼ� ����])�N�A���a�����%U�t�fE�K,;���bnu�(� .���8*����t�}v�ۍ��l�i�����+HY�}E2�P���� �����Plt��`^Ue��1�D�צ�2�w�����{or p�X\���c�3�`����>)�p��|��I�c���X>m��>���� ��p1w�����o4�k47���1�n�{E���/���{�l�;pmѻ �@��2��/���˸Ͷ>�	|���G���k��/F��K�Ao�Mn7�>{�[�T����gp6�-bєY���s��4����{T~G��b�5Q24l�����y��n�:^&�TSy���5�]���
�D��3�������~��/�2)w�Īd=:)ɜ<~�r6V��g��[�X�	���F	�f�,CQ�}B�����I:��_�(��GX.,�"� �c�ͮ�K8��-pJB>�*Gu�˂�O�n��+o������Ȗ��D�
'P�J�g��+�l���˜(6)��7|f��.-Jy�f}p׬K���ܰ(�ɛ����\i��ϐ2N	D�[�;���| w��f���ցT&43���3UӚ-��NϳVv���t`�e��r�7�3"�ŵ�߭�q+��r���~{��@���E��ڽ��%y���?�ӳ��b(#,~�_&��>�ɻ�;�$��>j{ȦJ�-C�[[��b���yۢ��"��v��K-P34�������l��(2Az�7@|}J���Q Eq`�Sߐl�a
H?�<�:v��e���٨ݮ|����\������u!t<D�5n����Ξ\\���ύ�h4-;¥o�F�EV��e�S�U P��X.����RlZ[*=�m%0�N�N�J�	]�9f��$#���� ��|�Ah�6o=�?�ύxv��Z(Sa�-����-/VU�d�~�����ɸ�0Y֐8��CU.�ε^��^�:z<����Y9O�e���p��8z]����=®�HffO$H��W	p\%�&�Z���q��e(�<�����2"<:;�ta�+;YkKl���G_�Mǈb3hɽ������'��#%$9�r�F�`���~���4�C䠯��XmD*S|����kկ�v��X,��;Xl���H|�����F���`@ˁ��ӽ��޻��#	%,��t����m�����gu�V��xJ'���]��8�b���;�[&5'�m��g����Dd�����^���h���v���67�y/��]�1�dZ��$0�zn�`#r.쁼�G���/a�

/�4sy������H�.�E�i�Q�N=I�};Ls� =�i!!��w`}�v�"��
�qȁx/��$*�;ů5��UP�Z��J�}��S�׷PK22q�oӀ3'&�2���5�ѷ��2��l�ݵ��h�ί3�5�F��a�}Gס��d���2N��?7U;N	��N��x9Y�g�x<=�]�0�p-���⁖-�JpV�xO	N^?A�:�q���E�m��P~���KV�BP�H�{�������G p����Y5ed��_G�b)۝.4(i����S\}@�4t����H��N��k�sؠ��;&
/Q%���3"?L@l��]���M6�2��&EM��]�>���~˃�Z��yN�+l�|��D�k?-N���j�<~9�E��M�i ��NEr�#l�ߚK�]sӋ��uk�2���|��oo����X`�X�iIS@�Lo��(����-�E��Z�1��3��u�
����ñ�[��Q� f _^�?���⹯�P's�-e=����jJ�ǆ�?�p��<+?w�9D��#!�׍�U��ԟ�A��b��x�|�p|G��[G�N�靇��H���|���-���Z������#�3�ӍM}o��S$��n}|^p��! h[p��k�1;b���u����=0s�7���@���<���j�x�#����8x��I��K���(��@-��>��i��{�bS��(���`Xq�����M\_¨ND��)�O�����_Id*.���b����Ӛ�j��N�}p���?��גu>K? 0����)i!o+�&
����o�	����>Ҳ>1��V�S:f�z�e�|9h�%h���[��eM>�j�Lŉ������I%�� �p���I ��t.��.����*.���ax<�cƱ�tN���$-�ߏ�e��a�Vdqi'Q��u�j��Em��zsi�z>�,�y�}�шKJ��o>����܂.k:��v	���x�@���5������+��:	x
��&	�?)%�o_~�1'�g���qj��aA[ȆZ���c��C<�·j��%�Ó��a ��EF
���2T��� �*�㜥�̛�.)��>k�vߙ��tY2Ay����B�Ӯs��_���N���Ō��@(��vx���Yjk�G&����9u�Mش�o�Ey�!2��� |�7m�_�ǟc�$eCKr�I���ҍOE�n��1��W�MN���rEO2�d��+v�/H�}��u2և�a�]�G�r3Q}���6�B�&�,�'6��
ل,�;Rؔ����O)�>&�Mς��� �z�F\́�Q��Q>b�]�
KpG�W^p��a0�O��4���Zw��+�V�W[j���p��@���Z��,�]���D�Z����T����U�%JFF�L5����E����{�{'و޿qR!��p���_
[SǷ�7�pR�����qF��]�5��)#x*�c?�-�PZ���V;yMfx�^���4���'���\ebX�M�C/��q�ݝT����_-S͞:�&Gpt4#1�ީ���Zgo�'>�~K*6��+����s7�?&��5~���;K�����o��n�@Ҳ��20�(��f$ �+���FZ��{�X���޸+���1)��$z����������{���S��@���=�rtቋ̓ �GU�B��Ųa��5٦�����#�g|���ep�w�;=�|�?'^�G�{�,ۑ�;myܜ8�{���)��p�%[�d@l��ؐ�c�IC`}�LM��Zx��ϙK��7Pa��z�H�󪫢D[����e:L@}?6����&"��j����CO����)��p�yfY�wl��0k簿��#a��rM�̿f1 �G��k�U.D*�<;�!��c{j�-�3T����VqɟÞ��+(�Q�E�Z��`}[�^C���}�X����v.��EͲ���,����f�Q�}Gg�?an2.���D��B^�lP��slx��v=@����`��1ŉ ����g��zG���U���j4�H}~���V'�_@�c��	��H�s�.oN�n��2dײU1k�yA��$A��W������_��8$z߱�����^�x�	��>m��b9��:�,��tF�ߔ�M�۔�tIT��������]��G��>b�G��^nxd���X���F����U�F�EC@%�|�Yn��ƒ��;���� ��G�3;��~[��.7������w��\������ҳX�ۛtQ�閿�x�:{ok/Ū��}�TH���4�~_��ل��r�?g��(}��O�L1�t~i��kb5Z����]g�����*�F25m%5�ͭ-/1}�
 i�A�#�����*j��^�i e��"\t���&V-b��䃦�m��ZؕZ�����؋�q���bp���Q�N�zs�����G�,�|�R�I��`�va�� ;j�W@�kR^�թl�הP�Rh]�^��H���=�r,�謻��3!�-��J�e<4C��`�w�|�*2V�������p����Ҟ{���'�`#�����~gٙ��1R"�:YY�G�2�l:��.���J[����z�"���՛
��i��Mx������=�<���[-WFhC�D���EG�+���<�\��fT����6�$�NO���Z޸)$��`NJ�i�5ϭT2�������}����ȡ(�f�Ȗ�RVn�@x}$D{�Y7$	5�?�̙��rC�o�~:����N�eQ��=4���T�ı=O��>���@�x d/�B��B�g��5-,�Ǽ��g�F��D왳5c�e��͒����6{[B�h��uX] )�6a$�qݒ��g.�V���~�J�uk}��T�6v �zk0wgf�_���f�5�k���1ة��s�4FX[�J�����6η+���J�~w�v��׃�rͱ��4�.Z\�Tv��8�u��
LY�V$��c����$�?�]y��0>�y�o��`�L�̆ä��p����\�|D�Gp-��q�.د[�Y�����R��Ci+�h��9�<K���Rv�����Hm6����d�^)~O�-�T��)�!�Ë�[�ʖ�ݧ����fGR���\.G:��23��A�t謔`e!)��2�#1�çl�����?e��%���ۇ��{���DMd�Bm�m��T�~^[V��Nh��4��o��7��Gh�[��͙�u��Ƭ/�?�[qL�4rH.�82����tg��g��,�1���̟�`�~�y)bb�+v��>얤��W����j[«vݦ���cSR�d�P���F�C���/�䟤�'�o����h�j'�Xz>W��^�z$^�QK��z�M�7��P��۠��jbYv���CG��ؠ����߯x���t9�����Š���������F7 <�{�\S�:�y��lˢ]H����C�/�l���7E�.��KYB�VD.�L��#�6@�� �?�Qlݾ?Wa��U{���R�i�ʅ��N�u�Ʀ$|Ɲ��0��eg9�0��)�j�]��f��~�zN�UQ��!�ha�N�;�"���1\���i/%?�{� ]F�&�KJXI[kz���ht���
G���T��+6���F�1�{�p��*\��'X�ŗ�<7YE�r�?�IU�����+l$6��.'v����&@�1AT�����UN^e�U��?����/n�w���^��ڷ?���8��P�C�ҟ���k�l�b|E�?���HW�"�z�`�mzd����c{ǩ�Gח�C���Ouӭ�����H�5�XۨlE��"Fd�1v�+�RY� B�H����,��%{�:�ƾ��9t}����^��2�s��,���<��+
�R�s3P�%����a|ޗ�5�������E��'2�x֙I<���\�=`Y�lҽ��?`�� �ď�R�"o�C�T���2s���ԩ�{�Y9��d�U'R|B8��;cm� .B�q���|M����{���.^љo^eKỆ�v|O���=Y�n{Cׂ�����B�� e����Gqݸ}פ��_O�
��]�v(/?�gO��J&`�*>Bϐ�F��T�o�3��~���E31gi��O�<l��;���.���m}
�V����u��(���%5�]f�?/� 78O�6i�'�Jc�^�Y ׸�a�q'��n��;�&C_a�9��{��[�8t��]-
�Σ�V�]��� %_��Kd��/<����a�mf��M�q�s8R��b]�:2Q�'��Jj[b��Fiv_�����Kgmt�9&����>��H�:����׏�Z�`�����v��aveh����2�7�X�Q�?E�z�H�Nͳ3�f����	A)ʉ��Y�<���� |բ���1���܈Ѝ�]_�oO�~�kGT����!=m��,nz�b�y-��������"���,�G^}�l��@dǂ	��x(2�5����/�'��=P��<W�� )u@1�����$�Ҟ��fJ!����zɹ���শY����Ţ��7jL30�P�V@�������KE���P�����W��1G�y@�R�\2�l��}���1��H,��X�<Jd�#�]��FXY_�߆p��4����K�6O�su�!�؆��5C����*>�t#��}�����Z��Li,1�4/�W���،��!������*����ZP�rք�o�q��J�������<�u@qJ�doS��b�Kz1�(�������9���L�(�����X�m~�6��t�ϴ@bn������[!���7�z ����4�$�I--����o]ѸbO����}�����E�>�9 ��I���sI�V������n�@;�Uvh"���J�Q5G���fg4W$N���̪q�`�M�7-�/!|Iz�&�w̔���� �ݕ�B�h�s(��t���j�����1�V���W�^��7tγ�����r-M@��]��c{3EK���\��AS���;F|L\�Q�Ŭ�V''�?���wúU�;x[�AC����C��7(����L	ζ���Ϧ��g���F�m���]N��4Y��@C��V�굎c��V�8��U�wP<j�����(��1eឈ�%�El�
�d��W��f/C¦�8�* �FJ�l*i�?e�x��t�P�`�MUh�] �B�Z1=&p��8�:y�ڦ����ʩq��7B}��W�cݦ��|$���x�D��?u~Q�����i7��_}����=������	频6�����K>bb���ʽ`nT��?�*@��3d�lS�X b��<�:@0_��a��T���j?|���WMӂ������1 �lT��a�'@P��jH3��ܪV�&��*��?�����?��	�ץP��c�pԠͣ�l�惢��z ������ީ͝ȓ�RX�@6����?Y���wh �U��ҭ���
����r��Ƶ
�6 ��Q,�L�w]�@�W"«́�q�_R���!�&&�a7uc��4f�,��?��۾sӾ���EE��4��2v��[`��E�\�|~v:nSP!�A�X����/{W�o�Aj�ᠲ��f�U���n�o��n�qvmv����8��si��"O�������or�#P{wI�Q����&#euU���/Eټ����qX܌����-�&&����l�w;>f N��k�Y�r��;��O���?>�~�l����p��߮�`�������,S\�X�Hqs�F�<�/#{7#z�y.H�f~���Ȕ{�¶|1z�ĝ�!�o���0�ߵ� O�Q��������y6=5�����N�]-���Y+���N��͔�:�ɡ��ő�r�Ij{�2u�������P(~�]4�.߬��C�~�	�Eiدh�d�a��S�^�vSsY�d$�������!��Kt ��$�G�l�U~�ґ!fa+$kǬ�r�U�3K�3h��\���YE���%��F�U{������T�yT���uG�c�O867[VE$�<q`V��t�5wh�j{���s�C��V� ��<���5�H�q����=> �F �K0Ӹ(��{Zl��V|�򳚿�ΞKr�H����!�nIͺ�9Q���꺢A�3�.�ioь)9$��u&�K,##u6.DܦH�!2��l����'�,��4p����	Ǹ�k�[u/fZu�X��%ǂ��ך�,����+�Qeu
cK�{�-�|e`�Ň\��&ĻZY	l����rʉL�(��c�3�uѝ���Y�hu�)�O��9����>>����YV���C�o�Yt<Q��{�ۑo�|+�%	�ۈ�e�[k�.��g� VF����ps)X�0��0�!�)Ƨ} ����ɥ����n0<4~_%��Ė�Z���e�I{�@�P=/ʙV4u�`���2D���j�k\O�vr���G�`Μfx��f��1>麄��ba��6���U�^b �s����0�)bJ��0Q�\��fK��[�3l���c�?҅�zU{����N��'ׂ"�Ө��5!�E�w�T���c�P4�j���י��ڙ�v,�$����
d�Ȑ���-7��*X�}���#ISnY;F�t!�:�uX/gj��Y~E�Z�3�@C2�A���I�i�����f�}�@�x�<_�*^���4��]�O�/��;ǵxˉr��A��u+�[z-�i��� ������[�H�rZ誥�勱�Y&��aOm�s��-�*���Nɴ�N1GO>�´��h�]�sD�ݏ�e��$�#_v�O)�9߾x�AD<[��xa�1j_Q)�[C#uG@[���	�J����x}����(�w��t��y����"�n:?L}1��*�/�%_t�*>�������Cl�ۖ��#ᑱyl�vYO��瞸���>�����nT������P~��L���n=6�
�E�Ak%�P]��0,4��>�.��mBw�*�0���An��D�o���Kꉅ�/��n��@!��� �M�������6���P�n����bÒ��+H��k
愖6�@�ﮡ2P��~����E��\L�Z۹#���C�v�5My�_��Z�ly�Fij����~�{�������:)��N����=!���6M��@���{����)���J��h��ZW��YT�@��������=U�%ҫi���#�M�Gv�āS�2�ߥS[�u2f��I��y�#]�{)��c������Vc�LR`�Ò:���ӗ˾� dS�.��;��0���� T�w����r ���󶭗_��\[���7c23��Ҝ�;�L�)�k�f�V��Ut!A��	����d���y��-܀�r#&2`�����(�e��+Q�٪�0�pz����k���������R�o�BvR�-��]#;
b�"H�\zK�>�s5H��hm.t���+�#.����#���&�_�ڹ7� �6���</���a�A�3S�%�����h1�vG������"z���\v���&nQ�$1�O�C�+�{2��^9#��1q-%2D"#�o#x^4m�5��R����\����9��^l���������J�=x��X>��No��wʁn\�Ǚ�٧�d��YGw��i":��+���,QW��`���׵����0j�,27M����2�ب��������� f٣У7��[/��V��j�I���ad���.ZM��E�K� ���7j�C�J^&�ܠ�Uq��>�
�y)�Z¾��5�\]� ��A��;M6��B�zB�#�c��������
��	�W�(�Q�S}��ޅ�u�oS�X=��q��F4 "���֋�Bø���ƺP��`C���ע����S��C���H�� X��0��ר/�x�J �8���Z�J�wi�BWH�ҙ��'�)�-�]r��1�Y,~�.6�j0����	��i�|�v�ׇ�hu�k�`?�j|��)���!'��v�{@���hF_��a��1)V��Ҩ+��R�d�[zn@i E���g@Ͼ���&��]g�EV�O%����b�a��|�/l�|#ׄ?H�$^�q�]�S�n���k)U����ʶD�#�O�}���sڿ8"mQ�U��)����g��9�����ٶz{���|�H8Lp;/��(:�Bj�K�(<d]����<�NՏ�OT���O�9�Z�e���ōQ΃Q@�7�\�b̎�C?7��g_]�+�U>	�x��F(��%�Ʃ21۱ �����(@Oy4�v����.�m��%�n��B��/�- T�ؐ���n�|7V�eu�zl*����-NO�=��V^wA:�a;h���_�5�=�N�у<�t޾��aP��^���qx�"�(���p����;���5����/���LY�e�+�^2��A�v�qF��K/~`֎:4Lb�q��,�>' -fk���ҭ]�F���w��[5&��[+��[�Q�Ɯ�Q�W�>���up��m݂�?�4d��l=W�7�K��K�&�e `�Vф��0o��@o1��P���"D{9ɀ�%��|���/m�|)m�ϠAP`=ߢ�J��'�և�j̤/[[`��=s�E<b�@W=�  �`�O^^�ow�w�匀�a%��%ƿ;{?���}��ftz�}�6�-��_��l�<
��z��H�+����'E���%R>p�+�QLR_@w�{ydZ-[#�ю��1�Id�`�����!�z��:@=�C�Ô��/s��B@�,X��a+?�VcGx,kC tX(B��r��}���<�i����f��5*�����bG��থ�R���%�fn���]�L�y�)@��rO���5"Ѩ�n:y�2sp�a������=�Α#,�^y��o-!2�dx�~Z�b9t�i��	�n��,���QJKu����o��L_q]v��P]��H���\^p]Zj�Yw�>^�%F[�X�hm�jjy�6�2~K。B���?/��t��n>�ˋ�j&��D;�e@�őW���
�nH\�����x�e����E�Y���1Y���E�%�5�jO�*����cQrs�W)���*}��'��a�;1R����0nY������ L�V�C@����m�'�{	�][K��v$��EUS7*m-h�&p?? N��q`�X����r0����)A!��m�g`�D�I��EZLk�_���8�ne��:Z>�1�T�7�6ʁ���D�JO�'[q�����Vsܼm��R"^z+z�����wP���ԯ K��b����@v�(d��.O]���HKe����F:ri�$����gIuN���c	�sȱ.B/G���ֹ�b��E<b�"�y�q�>"�������l�!��0�"z�:*k<�⎵-�!��r��T��86�YA `],���Ԟ�=�krJ�ΓNKCN�O�5���~�(��0��|��?ΘNխ@�����D;�$1�'��(,�������tv �:�����AD2KS��a�o&�m�yAIZʽ����_�X�@���0`=7n��Y!VP�b�t^_b~������]�:���;�j����0��*[{K�\�؂*ɄI��y���Pz[j`&��/ �Z�>Q��:�����Uzi%�,Β�
�Ӛ�0�8�p
F5�ɟ�C������;�[�=���>JS����.�������p):�šxW�%�m�y��5����#�L����8壭Ν��s{!���7����	�'dҎ2S�r��;��8v�N�:�!�S['2q�.Ad�$%P�pat��B��O[��ڠ 	c �;9�' ^�-Yn��X��"�[���|����؆C1��4�ap�Q��c�pG���8�18~��0��k�T�$A����ƩD_�0�}N���QOiJ��aG%*�f25=K�z;�,�{~�O$+=A�-H̍�D�����0ծ�|!|I =>�������*Y>�,�\��*�_���H�� ��S�V@�,t�����G�೐�P(%f�V���&@���?�Af����s��'�-��>��<�����@���筑�TR���%2�7z�kV1�F��`q���U[�]�d���2稧8�����5�x��YbL�9j��:Xw�>���:�gC���;X�bz�Ji,�[/	�j��z�~�mP�{�n>8Ѻ����qs��+m
��cY�������v�o��Rz9����l�pXL�Q��$�Ey'�o�#���6�A��r��K8Pn�=���O	���Rҍ��=G��7�CUr?�}�;��F���"���`mF���Jp�6oI�/��T�Nʅ�;�!�g���l��F� _؇{��������C��q�����/��08]d��d��lx���\�X���^!�	��u)p�ov\&nQ'[��:��ՙ)��ؚ%	� �݃R<��e%˟��DnT�I�9�-E���ǘ���6ڈp��$t� �������,\D���rf��f�c�)u��~����� (l��A!!�U���5�8��]����)+*@4���'���t�,շU���l[���'��RNW������B�����5��
_�����0}�(�N�=-{ �߾�J�e�t���c�ۨ���B"p$�.'GD�#�� ��B�4\F�I�M�������-�Ϧ�x�q.�; ��tނ�q����
��Nd�NR���!M��pC㡛��x�Lh�T�.��g��j�, �åaċ/H.����&�Hq�&�%2��1�(�$�o`i#�ka�/����\n��MeA��}@��ߍB	�IaQ%����Y��$U�xxE4�ӣc�`�#��吖[�Ǝ���w�P�q�-n)Kr@9�@P]{t�ZGƓ+�^N���A�:cj��U�]����9:����8�c
�NC�{�09�v��y,�a�N �6��y���J��k,q`���r����w�̜��� ���V��\��S0��BlC"���ܟiy�0e��j��xO��c忶Nۿ|F
�
X`$�j%�P+��]��� Hh��?��5��t����A�֌:��}�D�S�*ˀF�t���h��w��5i��4*�	�g?�
Ȭ.�����r�HC��T���g�佾m'`
!�
@�q�`��N��F�6��G�I��L^���t��$�GE���9��]���܉Y�à����#���ս!*KHW�>��q��q��s�{B��KɎs))�3-�@��@�]<�Pl��҄^�x� @�{���<xd3r�ۖ���ua���!��Q5b &�(��W�>�{��k�h?�*u���l��( �Q�[�~ƒ&�����X�'���_�)ݥ��z� ����	�,�f��[��=Ǥ�������M?�����>pC�?|�L�JRLJ͑�{3S�Ѣiw��h���ݩ��sL����`e��Q��,tv�m�a�H�#����l����d���~k-�]ܘcdM86U �X�T���3 J�p&�ŭ��⨿�T(+���v:�k����
)�rN�o�+g��\j��>���x�/�A3@��ُ��o�^�� �~УB]��g�y_�`��1�}���kk%ت����s�ioC����� clImk3�!3[ ��v�V�� ����c���e�'u�c2 �e-�"ϼ�yb���a	Y���
4����Y�]�KI"���5S��{�ޞ�Z���M�ɹ4���)�˱�f�Z�499�:�w�6���~7��:�M��
�:P�ڵkN?yǧڎ�5��Q4E��ʐ�
��	����.i���N�?
Z���6�9�mp��qn�����\1����Wf�in��=�ɾ�̙�f���_�>��D� �p���z`���&H=�3^|&�/b߶U(��%/uJ�Vj=��K|t����g����N����5���ь�[ַ&�Bބ�%��HJϸX+�Ho��?%,C��T�v�������li
f֌�:���9�e���u+b�����#�,[������X,W��"�����UI0���<�����񝬎��ʇ7niG�s8,}[��3I�K2�>bu|�������H,bS�����1��N�_�wu6������R1:0�擎���I,6nm�j:@���OWyS�a�/tI-��?���G�����~��b./p��jѢ&g���ڧ���/��G��+��������ic���8��1|��y���|��o�[R%�<r^�����7Is%��QGjR��'/tl���=�
o̩+���"��ߓB2T�r��Xf<���Ыs�,i�hA,�X�$�I��b�F��z�yQ�7Q͚A2���^�n����I �-����>a��y>�"Mܕrs�Z�)�n5?[k�Ou��y���Ē�.�n���_�&0�n��g?oN���Ƥ��s��`�/Rz�PBb�	�֌��QL�����>���k���Ba�s�N~��gK-�Ĭ��: ������ �9���0����$��:�&#����e�G�;�=ײ�q���7�PCz ����>u���LSc��Ϙ��,L���׼�~��i���33Q�Νn.%`.�_S�)Q�/��C	ؘO��
���ts-�����M��S�
�ۧ��Ko�����l��\<\J#��+�tYA�۞�O�����!����� �?X~&M��N�э\�vw�q�8�˷ޛ~�=(�\K7n�7W�/����Y�.����LQ�7�� 
��s	�wY�� ���d�J��s��d����ş��+��j�/��%ej���\[�i�c���΃���	9 ?�JN�<Ȗ5��������/#F����N��Xj�M�B���In�u�<d�L������}W�G�#��r����|�vo��v�����N22v�[�U��ݶ`�ӭ�$�l>)�V�}T��^��2�9�}���7�L�:�G�!��h'
ʍ��+~�����ɦ�X����v5����
�������<�6��8o�Ea���V�@��m��l��S�e���n�s�3({��+*R��ca�u���.]$��E]��{6��Ǘ�Tu�j���Sၲd�`��*v����8(00��Gk����r�7�En��Qх��@t�5e���q�>;ܜ�@	2�x�l�(y���v�C쓹:8��U[�`�z^��	C���m���.�Z��C��l�l»�P���P���rj��'D�|k����˫RsZ|�`5Z��ocP���Jb��e���2��dޜN�����`@�H�f���l��t�}��҈�C�kES��Ԣ�ܴ�o�������[�M�|2�*��F�r�{��Ƅ
������b���:�� _�/���me<�x�v> ���_(!�v��=��} K8U�Oc�g<�\�����p%�o]��%���P��)A|i@���01����܎�?�����?[����:��!!���,:|��K vݼ��o<��$�5Q3�5�`��23j�}���,u�S��0��,�[�i5��xeߓ�c�i` ��z�����.T�sA�a���Kκ�ϳ.��k ��7�C`"q/�=�Q���|�	L��T��\� �]���D�Y4R[_h֚w������Ê|G���w��~1Cٯ��!������I�5�PV�䣚Oȶ� ��'dW����H�T?��o��"C$��A�Ŏr�;��y�՚ݺ(��)L�sJy��~�N xԡ%ni�'A(���\[�[_��9��`�#��������b��pF<���0i[;h%c33�|.�������C\m�A9��]Z�V��k�U�%��^Bl�$���ά0'�(ڃ��Ր�&���G�j�j�iq�l��#%<��TE��Q�k�$�6�P��ރ��S���.;�7�j��s0�޽��#�p�2.J�
��Y�p�\9圶:��m�D)�(A	�)��������iU�C�������qcՌ��~��#_k�)�!��U���J������|�-Z��/MC��1���$��.��c�����U{�j���T{kV�L�l啲�����_���^���Dzqױ����M��U�� �(�T
عm	��Lq��5��ĵ�V��x��[!�>�FJ��l
6�ww�9������rH����4�:&=�{[@��?�͚��g��#���ȋs^u�F�}�络ʾԙ��H�/s�*�ĭ�?Uڻ��\z^D+|Kmt-�/ҏ��,�|���M��!HD\�Kzs:M�"��{��?'O��6x��)�<�J���_�����B���+�����;&7��r��z���J���P�m3�&���-o� RQ�+���}l ^����8H� ��3f�۟v���m�0Ф�ت�s�[����8�b��+A��q���kGH�?��'�;Q�d]���3Diۋ5b�$wmE��p�	Ţ�C�d������J@T���g��)nRS5�%�H�ca�j>�<�kڬ`ʼ -
�����R�ih�r:#�X|z�s�Eϯ�ks�T�� �L~M�?!��V�z3�b����A��s��1���*��.����QRF�>p,5�]���4B��C�e����L��%=���SX~�`￮p�q��#��B�p�X�p���e���v��X���H4���]��UX��NWII3�,����a�(�w�?)�|��W���]�fR|�`8� #���w����@���%=�O|�'���IXa����_��k�퉀 >�f`��}z��`j�5ت{��:$<b�gmM)x~������շʣ����Ҧ�� �>(m6��R0����2gF3��rT�`�ބ]���yO�o4�o�`�K"#+Y�� E|p�;L��C�ԋ9�/5 �r/���,�P?Y?�����3mv���i3a�O;&7��5����� �><]ѯ��3��{g�?ڂ�rY�|e<�"�s�Sk���c�$5��Px�Qx-r�s���,��[����-:�z���ܷ�M�P�\W����aF��t�-Y�z�t|��_8<KuS��ި@�?|�N�2�����G%��M�'�@�keڛ�0���k �`��+l�P6n�^ml��ޑ=�%n?Y���ث��a�IJ���Q��pinUK�Z�qG�p�Y�~@�|���Fƥ��p�?[��}��n:ѵ����~�����75���<��Uh����<�����;^y��?�C����.N���t��� ި�LI �������_��:΍��|�S0�s��	3�C�+��W�?$���}��k�����gO����9Ɖ0�+���W���頿s�l_,����`Ԡ�xr��Y�C+���_��]�R36 s���PnY��(K�%۵�EeD>��!��Z�N|k'��D��܎�����~�X�%�ih��\������������	}�Q ���߮(�nb�wX	o�R�g;�i���- �`�d� ���<7��(d+"OD	���=����>�Tj �#�!��ҭFf���!W@���'~�_&�w_ؓ���ьp߈7JlC��G O��jb����À`���kc�bp���rԍ��������@� �~e���݂#g|5����w���|���L������R�썃�ġ���j��w���a;��TO��x�]�S���|����%}Zf��T@{Ǐ��f��vۘu��wR����
o]�q9�y:�f(�eb��+J6��N��9��(7M�(4�������?�0�H@j��`��\�~��{K!Z�3�v������a�]�hG�[��ɔW7_�
5�4���"�q�*����p��=���ʝ��ͧ�������w��%ɩ��϶o���ޮ�0Dv�8�����;�~o��_?۵���
�u6���n��<|�K��8���O���~o�E���xq���-�I9��Ϟ>�?&.�&�(����Л_���R���ߖ��?FeĿ_[�j����7W�����n�U�����/���,�?^��{�B�I܏�S�é�7�7�<;@#8��]�mAw����&c��n�.�Υp65���e�j���8(m��Z=��dr��>!Rz��R{;Nz�E�vԳ�ݶl`lu.
#j��b�{pD�l���K$@���/:���@3C%V���,��O�f���hضD��R�u�F���c�~��Rp��[�Z�~�� �{�2G3�W�����?Wa8N�V����y��X�B@@�����m��=[O;SFbT�u��lI �4f�Y�Mp����N:�,��赖.��� *'��2\7��l�m�1	��UK���tb�"�Fˡ��BB8�|�\.+��i���Z�K�w>u(M+8g H����'�7�X[�4���'O���	���E@xk��&�����3[g��3Ϩ��N����
�WLMM)�Q(�p+"g����;j�?ῼ���"��ө�ۧzk�~jw�P�3��E���&�뤥o����^��o��U����3xAA��;�;�o�V>K��|k0pӀ�"<����z١��e݌�'.BZ��n��0)�(VE�tq�˔_�?�p� �Lm��> ;?#ݐc�G9�B�]����xu��G��rM�����|o����˓+N/ޒ%��YgYK~�B��rm�����#o�p|��H�0��I_/�r�|�[������/�)g�v�ʫ,_���&J��܈Z�ﵑ>g�����aP%X�\���g\#��ǈoE���f5|�G�|t�kß��������ԕ�?��+�����eV-^C�V��5�^��s�
�'4S�mG�����^����j�k�k��3tf�
�в�+��meQl��`��IPmZ򬘈���^Y<�\Q�Cm��m��i���"��=�աD�$'�JY/ᩉ+�"���2�3g�U(n�0Rn���d�Ę!al���G��%���e�lr��q�{q�[kSk�`K˦�q�%'+v�Yӎ��T��eտ�k���uo�y�1�E�	��`V<q+*��LY�W�U�-�w0+ˢ׻�_��i�r��=	��堪��v���IgN3�L�����u�6'���=X};�k,�6[�{�ᔊo�r��(Kc�<�a5�Jl�B]ɐP��L46t�VN,P����7ntE+�/���X�\��KL�Y�-lO�lo!(G剪�щ{Fzz�����W����bt秕��q3��
ǰ��#z�����.��9���s���k���(M���޾)�Y�GV�Yֽ:��:��`�m}�\��_�/��X��	�[�����\��	sE"�[�"v4D�ؤ[�:����i����}�]MX�3��Pu\����{Z��:P��ԫ��qy�jtU&�';JZ�se��!������P�`U��wY.���c�
n;�,Ώ{t�	���F��~��`����#)Ïݵ_�f]�L^@�`�l�)�C�u��}"��u`ս}'}_(����sjK���8mI�ଷ0bיhs�v�Ѩ�ĉ��
i=���a�)�.��Q��M�Q��?���.lS�C���`���}�	�Q�y��?�՜YiĀzE�W��뿔�I��L�����jR��}#	�-Js:I��"��Mx��t;h㶡\(x�5Y���jz�=�3E+M�uE��'x������w�E���R���8�/�i�Q.�ϭ:�S=#\�P�������?Ҿ�(c#�L(���@[�^	a�S�Zj�#��;���+>���ڽ��:K�9�}w���a`��	�T�%iz��[@�*�7rC����dʩ��8�x	��@�-�0�9���y�������-��q��QOԖ��d�25�a�k�2���k[��3�u��߯ R��$��7N���r����:�d����g�9���
��B�P�|����f���Z&p[��G�X����z��Њ���������.j��c�\�"�i�!M͇���e�u����0�;��S��ZG�,�-a��2�'����Y�B��Aja�.����Jd��cF,����� �`����[x�ģ/��%�iHD��I���f�nr�(~�&G7�f��̏8�a��&�{?b�Nc����l��F�\�NA^O$����ܠUCj�p�s��l+r�CR=�>���;@����ʆR�� Y{e�
p+���é�g��5i���O�k�j<�@*wZ�_�_؁�R'Z
$!�3��a^a�����<�����f��EC�I��ı��$��FJw[$���sv$�:����'��-ֆ�}�h���ۅށZx���&p��n^��^^HS穿P�펠�Hj	�����̚�(䠏
<C���鍛�Ɗ��o"ѿ�gEE�u�E?g����)������В�ˀ2����1�"�����M)| i�Nuu;I��^@Ԣ�%��g#yS��� ��W1����c��@���B3CJ����">l���b�܎�	�N3I��G*8�鹮"G���(���%�L�f9����&�����ږ�8-SO��\β�vz��dQ��n����'^E�����qG6?p�Q��7&��K����*~�8#3CL:����B[��H�� �&���B�DW�醧��R��NͼK�	�݊ꑣ�����U�?2!��-�
ؼ5��13��Ē�Y�h��׹ˆ�R�]�0zy>QZf������n�&9���ϋ���s�W�{�+���/�L�����
�@�?���K���.�����T�9�8[ee��L�c꿓44*���s���(��W��q�~h�������V(zn�����K(z��Ϸ��n���1���6�oZTN7ko�Ũ���x���^V��^$���\ er�LLV��-M���؂��)����N��ˣEݰ�}�X^K��S����>�]lkכQ%/�>P�R��y���#X�
Q��!¥����a^��L�O�]�R����ǉt��Z���{*+��\����I���;���@_��~÷L�sja�����rV���X	q5w�o���=7�G/�:;i�3
��V���bg:��3~``��Xq ��\G�ݣ�wi6o�~~�}W�<ol��/\�]���=�E�0A�8��+�vs�b6�+ �6�V�uD�F4=��`�!�O���� ��z���}�;����PlA�m����]J��u2��~m-pVx�?b7D�֓��i�K�0i����XU]4��9�l6f�Vx�F��+o��C��/����eϽ(�E`ã�(Pl��mG?��q��x5�����iN�K�Tta�m ��Dk�O�܏V+~�3b]��|pxGH��s���--|�X��#�l��z��$��?��^��������3�UA��^�6ˑP�fO�ʹi�����TS���K�p���։Ȼ,���ϖBɢߥo����{�Ѥ�:O�i$��
u.e�Yc�� ��9�,'�8�oE��N�X̌�r�����J#M�B�qo�Q�5����^�뢑�#9� �J163S�۴�V��|��h�r�^:�3�����o�(�)�-ݔ۳����"��醠��B�L���k�3E�\B:�٥`�ag.����у�
�"a-���8ɟސ?i�*xhs�.�9�o��m�_�1��p�����qaC�{�>��3�z���m�6�t�S���1(��P�=M�2�zrb�g����pV����_��>��ͯ;���:���VvK	���L͗Ⱥ
i�Xز$Ix�vFrb5�@V���W�{}-��x*qJ��9�w[�lϱDFc�4Y3sv�ǖ�c�>�|����CRNb�{,�t.�#wO���)O"�z���e���3��Ux�no�ɟE�,���|�bA,�ه���2�< (/W�F��ɥQ^H��WH�.mA����,,����cuptMe�?�b:ޗ�STj6NzBj0�p[6��9J�us�-L3�`�=��8�q���q�P���g��+��{Fu ?l��ʜ���ǳeı[�>d%	�8�ܞ(|/�� ����T��c?������p�/�4�d��D���5�[��K�d9�`_�q�"p����N��)����]�1��Ϭ��~���C]'zC��c����
�E��`# �01���� ko����e�튁1��������!���;�G����}�(��d���r��*Ū�'�FEz����6�����m3������Yc���:����x�V��t����.��nd֙{�_���I�b�]��8*��0���0�bK0r�C��78�5o��O�0�`�)�Du!�Im)����&�W�1?�A�$�d6��x61q�ms��2�觢��ۧ��E&
3T�V��k=O͔���:K&z�W�(��Ӌ�Hg~(���$�� 8&�pc�����Ii<��o�%[�=�{���U�X>u��Pq�����d�#&�R�O�AN��_ ��!`��I��7^��o�TT��SPR��c1q��q�9M9Y�-ͪ7�U9Q�5�n�Ҩ��
��[�H5ɀ�u~�/�4�b:Τl��C37���< ��@���[d��Y�,s�j٩8�G <��$Uͷs�,O���<4�8�RT口'�:~ѷ�t�"J*���5�2Xlb�?777�M���,8���07l�z���l$��S�������Z�F�D׍�����'D��]��R�ȩ��U���x���%ĵR1?ZS׬&��8�M^U3�����k����f?YG�+��cOj��c�-�\T(�|�l�4���wA��JP~/-1��a8ޘ_�ѵ?��A콊�S�(��P4f�H �'��&W]?�D� �X�'�5
�D�*!:����]E��.�#Р��*���� �,�'��|^]n��噓
C�*.�p�u��x�V�?����hj=*l�Դ�G��ѵ��COz����?]�_�oV��%�g���i�n@m�Ԟ;G͌Z��V��εkJ��M8v Z�ɟܣT컧��c��_��Q0<mB��_�ZSQ֘�?���N
B����M H�7�` �C���wW_���R��	O�nK"R�;vp:
Ѩ�m����Y�<g�Fb��-���4����{D4�f�[>G�gRT�������v���uf(�Pi�ųc��6�[nT5W���J���}ц\��86�vīKD�O�7��QǣcD�E��ˈx{���3؊���4�sqHt|�36��B��Y8 9?�f��?m���:]�m�D�Q� i'�S\��]�?�~�hc墵L G��5��X�v�8۲>JCZ���d��~Yׯ��6�n&�,��qMG���1����2�RX��׎\J`y_t �� �p|�i�#`̲��8!p��*���Z��;�ʺ�c��\�_��1$�V��B�iV�����?�9�f���\0���ɜ'�,}ɲE"���_���L��D�ّ���K3S�DfH�⏊b�+����鐌U ���f��L�����N��N����u�O~x��ߣ��e0, ��y��[����v-		*��!�Jq57�e���B�o������6������n+�y��VItf��$��g����Oq��!�z�����{ͯ���@��*�6(�~�n�D�~r�����*�I�?�X�6�6�J$ �y\o�z.5SV��	=�f)ݦg�
���)����"�yIU9���A� V�cQ��UM�>�eI�NC>a��
����F!Ȟ��F�g��]m`S
=C��*���eQdZ�h���_�l�(<�7wΙ��Ű���P���1��C��\�}�m�:�u&2�+YȎ��VL	��Tw�����i݇�̻^-X=߁�;��7с����A=�#P#e�]��ȏ3dD�;#�ϙ��88'�|��?ϧ�:������Q���Bk{m�����D��y=Y���~��'2β�����Tcu��O�a��u�F�֡��mQ1f�(3�S���{G8T&μXx�!�H��si�X;r�q�d��S�w��>�z
��Q�Ԧ���85�Q�qj_Y��2����1�p�����w"�WȗˮOK=�'�w�+�Z�YN��rHݬ:���~���M&r�7�؍�?qP}�� �Y����J�y�Vf��fs��E��ݍ�%Y����T�?�����4����T�mUj$�ۗͮ�O'%ze�4d���v�ɞ�~^9+��ji�)He��>n��Y��u�xz�~���{�{�`�+%��m�7��?S�ô�I���tY9Q�_u�#�}�K���CZƟS����W�&���^X�,�����1e�-� }L�!�qt.�Ҟ�; ��/k��{oU�Ǎ)%T*��T�I{�$#�!ٲ�;Q��d)�}gȾ3e+�:��0���/�}F�������s�uuՙ9s�����|�s�}f_�q׼�S�^{u=�idL��Z�V^nn���Q�ִ⛯p34L+�?�k0�e�o3��THm���hgX96� g�w"���ﱱSkN�<��#�[�̡�{@ �q��?S�j��ƞ� � ]���7�N���eXJK#�gT���hJ}A��X���}?j �����2��{���l�Ŧ��-u\Y��b���Wʋ}�6;H$2˼6�{����N�Ujf��<�zU���N�'�\�ۑ� �	;���N��ϥ��|���\o4^Ƅf瘛^S�IW�ة��yIݙtޟ��F"��C8\��p(��/��B���>��L��y���;��n+�� �^C���F��j�����	���6+z�t�O�(cP)7��[����I5'0H��Cw��t�FGj�J��|�Q_@���.�{��q�R�� -�bg�WNJזI#߈�u�$>'K[��U��]��W>wJ���S�v���\�kǄ=�⥟�)@�C��[Sr�;w<G��j�*��I��z�D��L[��#�c�|�"������N��u\.�6�hc����:����kB�����9MT����1Y�iת�[+���v�����;�T#2}5����(f�����_����4�9��Y�]�����y%nߪkK�X�vpE���cH��hNi�Xe���s�d��`���a�z k5���� ���
�e�ǳ;;\���%��S��(�_�H|���	���Sͭ��:"�$�x�=�������E�;w�3��\*��]f\�����ajs������9��zck�l;�v�44�Ez+��<�4��f�:ڦ��t�ѳB??��i5�x��h`�*�V5�@t��������\a9Y|
����a�kDռ7�i�h�3ȖQ�L�"��p]���f���i
�z�C�e�ӫX164no7e��$|���[�9U �uv�C���U�O�.!�(���IK<��x۫��9X�#��`�w��J��cr@<�ӐXwK��K���z �Ռ'-����\Ҟ!Sϗ-X��UZ��g���Z�t.�]��$���'�e��rLI�9����Lj9�zy�E�c䴅I9b`d��d}��R�m����{�M:���v�-��/�h2F���F[x]^��N7"nv o���'��^��|�ҕ�#�4��o<�)�O��'nO�����M���q��ݽ��/�Z���^��{����s,�������R�Ʋ�� �k�����e�-��ˍ�j4'+�]O-,�;\����c�֎_��>�"p�;_���Z�u�g��N-.��7�����8+�
Y,�k���s�<8�yN.1�5�&8�j��ƀ��oY�62:�<I\,G����i�E5�
c^�����I��&�T�%L�Y��G�W��N��
�	�Vrh�<����z�J��.磔�0tK%���\�lE�0�K\7��'Z�]�ix'�mz��d
]h��!�N�%�PMC�9\��:��@qJF�׾�K�p���b�%Y�<�A1�}t����;��ҝ�����D�q�5i�մ�;�3zH���"�
�R�Y�iv��&�c/C�٣����-܄�Np�P�y�Y��B�L=$�!_L�T�v���Q1��\T4��G��sY�W["�,��Y��W=�� no����70�m��GO��k�2��3�^ǽU-�-�1~� �3��*�!;u�d�RG�)��FM��������6���Z����}����a�GB�&�,>��ӓxk׎�l���hY8q����(P�̼ ��Bی�egR093~�(&[��ekrZ7��}��d?�]�ه]/�g�9�Z�,Ʊs������i�
���A5�6���45#n���H������p�@��44��Q���'���L%=��˟��Ar�E���Ф��T���u��Єڢ�7J���[~P`R�X�ʺN��I�������?W`0�ſ}��}�a $�o�ԛ�����Q�豫������P_᫇��-��e�4�$U�n�Ӫ��pn�.�����h��9��6�0��JCv)m�?�@���;�	��o��%d���kwk.���̨Fg%�����qh���yR���1.%s�k||HK0�������Q�u�j14��YfoWz�r�f�����ۋՎehh��0�#A���y���\�R�ݣ�f�8��˷4w����C�'#�?�C��黌�c��O���֋���솵�<�����ku��-�F���z�0��_M�-6�&a��!�ͬՁ�&�Q�@6x�͙~�͛*h��$��u&����|������g�����g�CO	$���2�h�]2�<�t�qLA�!z�#}] L���O��tN큪"�w4��Rx׸*�Ё<���+<7�K�n��(:a堧	 \�מ9�i�lee�JM�:~��z#�Y���y��wOڛ�J{q���q���N�+��*�#A��^>���<�y�їkh���~m�~mx�-VMS(LGNS��gRTX�cLE�e$[60(���ݠWh�Q^Ն�-�ǃɦ����tM�����OAQ�2�v\8CZj��A�"=v�Y�u�����˜���~Sj�F�~� �գC�m�d����$3m��P#�M_ZB�2�>p�lW_�"�.�Q��7�0��wĄ<aON:����z[9�*�<F����m�ھ�$3L�*�U�B.i#���$~�h���6QͰę^�`(�[?�����A?��׸����-Il�]J�[�\�iXS-���}�JT�ڱ�FF`�R�$�\eѧ�欉dj����y�G�r��j�ߴ/��Ὦ\ ��B��$Djq��R@!��2+))9�r\[8̮�3�����(Cd��4�O�oB�9�`}�ϖ�t���JP��k�TO���_�l����������0����B��6���:7�׋v�'�sk[�������PߤZ�jp��]�3,��[E��Ї�Gg����x��&�j6k&T�QM�l�$U�V���Un�N�ΙE���o��=����"�������VX
��m��"w�th����۱0��Kw>`�0���GU��k�Q7c���4t�I�<�w0�԰�1��[E��W�h��F�����i�A���'��Lj����͡�s��Ù��Q���]e��[\����=�,o��-��IPb7�.�c9Uh}�)6�2��Y���sܮ�#�u�5*� �-�L�`ee�^P��m����}��V߆�8?�#��Z.�9L� 9)���R��JAc2^��
a-��"�`75RA#�ZCN�4���:� �=OS�"�F���Xښd�͍��`��g� �7J����r�:��OK�o�*I�Κ�y� �c<y���^ͦ�,Z<���*3�?n��/L��ɻ���e��:�`"�����V
�rˑ����*L��5Y�y$�ء�g�y>l^�4|w^���[�a�/��SM8��pV�ϻ`���4�B�8��t<x��j���0ZYhƿP�!�K��b�������(�;MZ�����)���w��2�w���4���]�r�}�I�\�톉���i~�	r)cyqڰ��g#r�|��(�������G���s�L�u*�� ��tFJ��b����J��}?4��^����#�Y}��Ι"��dW
'I�+.R~��"��̿ǜO���%sRwę�ǁڏ�RwyR;� �%u����W_�`�,�
PaZ�\���.�饢�� �LT�E����I���fJ���j��q���E�4[�_���U<�G8�A܊ۛW�@��I��<[�8���M�����|�~�K����Ly& �0-���-?�f�+�Y����9�Ff�[s���Ee=�o햧��:aD��,��B"�"�K,�F
�;<��xX��Dp��&�^�MS�;e���'��y�����A�8<]ֶ6��Cq�S4k�~�b{[85��U4�|��7�r<8t"5�	�Y\5N���l�n���@�]�o��!|L�#����z;D�-į h��Y�!���,�����n�٬�YH/Ú�F<@�)-0Hs"/eY�c���q.�����;�����H�Ռ�sc5�Ɍ�����c����<������|s�7�}�q#�'N�n�*���!�[�l�:&��ς�D����ܪ��j�Cgt�ڂ&&VZ���? c2�^��ոWl}/��Cdk��#�s�@�L�[��쾇Xb�q�.L�
���C��fʖ���Ѭ�"��|s͞V��peW�BwW�k�3U
�������[w�zO�N��_Vӳ�gEVf�A��>oٝ�K3X������g��D���:����� �7��}uw�,�ҧ<Ǵ<�qA|_Cڌ��N�������)L��Z��������C����4z�?ݓ;O.�0���lL�@���ή�ܨˇ5b�_쾶�-b�g3�?l��?0�&:������o�=��l�T�Ev:��;��;�	��*IV��TK?��֧z�7�*Y��B�ᦇ�AS*��0#�ZZ﹞�H4޲5T�d�� �ދ����O��<��,x]��6���~	3>���}?`���+?6Rua�K��)�?��?7�ߎs��"y���h�T>\=߁���8�i7i<��|�"��� �B����������~����V4�����s^&�AnX�Ț��R�0>�o�	�nV�%��P�Ȓ�,Ȧ�����$��8�c�g��d���J�+��z��W볚���,�GU�4-���,��z��I�����WK���6dO�^4�[J�l�{1	������W�$��o�e��[��n�.�z�ٙ��h�f��F|-8ۖڈ4J���������M���KP�=3�4~���N?f^���8�0I�wvψ�QY�$O.S�M��q��Z�K�K[w�K91ocM�����4���Tv�X�Z��;B����XA���3[ ���^�q{V/r|i����Y�\# 4-{V�bnU�a�O..��UԚ�t���:hVL"���i��!�P��Xǀ���1�SV�_W#Մ�K2���*�O�X���loY����eY��� +-���*؏���#�*�nϖT���g$�>��<h��C�/�\��YGg�P�-+��YY�s ���m�ӷ;� ~\?��~�	^ �7ESLa	[�s�~���/ڡh�ۮ9�Y�]��$ �Ύŧ��A�+���5�G]�P���"�qr��W\����>w]��Ȅ��#�*����/Pkv�/^��2v$�歝Z
��O"h�q�o5��J�$_��{�̈�s'���@v�����y1h�iɭ`~� ��t=���|hU=����<�[ֻD�K�'� W^>PS��+��l�xh�9C�vb)����T	mE Pscy6*.L}l���=���oq�ߝO;$�����P�c�������Hv+
OM?9�nj�c!�u�4U���Iʾ?�5�cêk�͢�m�dv}c�B^F�)�b�YE�=��&Y Ǫ�h;J��F<���� P���)e)�x4�4�e�Y����<��=9ʍ����U/)�y�1��K�P7���9��G������2��q\���<[h=,�־�D��kr�կu��xM]�5]��Ź'�Q��@�ڹ�[ ��o�㚛����P�Rz���/$��;4�p���2W�]Ci����@o�k�X��5�Pɝ��j�/[�2��o��,_�Z"�f�=l�����J��_�*h��è=v�+O,0���Q��c� 1/��:0X�eˣ��2�6�6�j7�s��^v�a tE����+��Ӥd+�4�i}�x���r~Ԧ2�\��-`l�Q��ve���@���[|G�/�K��� ww��u��
D|n�v�'�|t������ �Tx������p��i6�� }��k�ʢ�y���y�]����7ې�w����3G� �8̙�rR���BUE���Q `'�M����%j���W�Y���ym�����%��h�)u�L��ے�谝)TI�x��� ս���Di;3�`�O���f���� ���#��&������rZ�� Xj�<Фf�����
��Z�Xy��0�痓����Y����I	���1���r�^܃�pk@/R�_Wl�v������M�К��W���I���_i��yc�X�_�x�k7�Z����(h��&2@�-��.b�f��1n���:Q��@�����Ԩ��b뚃�����mC�wԶ�Y�:�b����s��a<V�.f+t��#:��3'�x s�,C1�RjH�'C��O@K1~.�*-��@����o}��v�;�ԛ ��ښ)bQ=��:� �r��*�y�䷛���J��l7vL�![��%��EO ��Oyet�	Y%�Og�5�\k-�<��2=9�Q��Q|�$I��)����^�&��qN��Y4���!�M�y����� �T�(�	���`'�l�邆�;\QZ��
z��a^عC����$Tc�ŕ�]�T�RB��ؠ���d�CzL1`_��Ӌ��A���GO}G��0�a��%G�gz�J��S��1@�Y�����oy,�⊢�R&UM:��gM�mQ�'n<�`�5F|��Ō�Yn�
hxꤤ��-���tl�մ <�=?���7!��1�ֺ6p���H{��R|�˕1�L�0wk�|'w�N�G�����5��沽 }�%f����'���?D�zxj�Y�|@�#�4�Tpz"�6DM��5�Z辅���B��j�3^.�~���G��5�h�
��w;Ў&.��i�eo�9P<�a��ſػF�^�K����r}ĉ���>G:
�Q�K��B5�i �Y���MÜ�W2�k�*c:FX���:��#��3a�yv{��H��_��5#��7e��$De���M�O��.v_�=��a-x2,)�D��M�4D5�������z���,��:
DWC��GRr�-�P�>rl��f�9xX��P����r��]�ـ�z ��VֈzT�����C��<���[�? #<�T�����VK����QX
E�@�]0�(�Z��'[MC7@)&d�Nww�t7\�$�wdK��j�d�~�g}���w5�"�cx���3�[�Ά�T��q<oÁ%�Q~,�c�1#-*%��3#���	�z��,�.|3B/�W~ѕ�6E�%C�Z�{	E�)�v��f��n{Aap8�&D��G�  -1�u\_�`��b�xP�^�6	�e|��0,�O�y
��_|�����x��0��<�b�.0�4�ZBҀ]/���j�ݵsj����l��T�T�_9�@ᓭE���4�pq�I�eXȂ'2�3�&0t�6>�:�\��5��B��$瞮8���'� ?z;��F��ڂ6A���
�S�DK|��+�fB�f}C�v��AW� �'�q��-��#$h3"Z�z��E@�W���O����x��6͸�Y����m������z���f�pec��&��Ł�f���9���V@�1 :��F{�[E|*>	�eh�8w9�	��X1t�' �N���TYoW�I�|�W&�-8�4�.�q�룠�����A]|�H_��C�y�5�^A�Aey������	rץ�~PV����ŀ-�Y������p�����('����B3��:`#T���c :A�ud�i����Aj�k���Z�dO|�}/@wJ�5�rHp�sa�=�#DBm��$X*O	v��ͥ��ޒY�$�{������@����֐�⏑*��1���^�1��	��CE���F m�\K����K�K^�G��)��i!̎ ��T��wX-���2n�~��H�y����\�����ez�S?��͎�V���;"1�
����D�p�H�d�nu���k�;r�	
���X%��4�J7ᢊ��R�m. �x�2b���x�^��H����ji�]���M�!�����t��QN ���a�O݀BU�1Y)�����!������:�����w��P�Y�'?�*-�pY����x(�v��DAf�.������nx����ݵB��q�]���4�&�~�/��߰�������<��1�#-A:�0t�@%i�  ,��� lњd�%�I�U��<Cy����)������S5;kc�z�����?QrsCϿ͗B{�#�Ɩ�J*���:i��#c^.�t���K��V��4I�-W�m@I��f2D>Tj'`�����a¥����	x@"`dxR�"dԓ�wg�a��F��15}ֱ[�;�e���7ӫ+�L� ��k�P Ym��>��:P���xoM�<�%U��zf�Z�>�9�+��]q��'��>R�ٺ�k=�ꬖ�f����j���Va�k�^,�L�@�=42�
���+_���hvoe>�Z��M[���:UD���1�
�����oЌJ�j<G����7� 2 �3��7Кɼ�&[\�6�_�SXC�($�$D���J �,�f͟��l�8�?�杨����z!-)�j�4�AB�	�=0|��$�F��V�����/i@=f�U�Ý���Co��*�2:QQ�|9�e�GK儊Ņs-X�L��UMb�����>�@�-}4m�I���JiA� ��b�cۉ�A�������5�Į����x�e�aa�����cN�˷�0蠟h�0L�:u����o(����N�n�uw���� D�D��;���<���R%��J4�!G�o~�}e��$ؠ�Lq$~�S]8�df
'un��Yy���e>�+�"*�m��wS��k1��Y ��^�����>�x�}���vj|^Y��N��*Vn�n�>�/ӧ�.�ngno%U���-)|���q_3om��/{x�[R�	s��U�6Z��J�a��.6~$���:[�\����"%z�`�������P鋖�����_9��9@k7ɝ=1�B+�$N��닥�h^���E�[`}�����ל�4�>cu[�:	�<;1R���$�^�M�D)mG�\ �yA��!�PeP��Б��@��T�S`VrƍZ�5[�\�4���h	��B�ĺ�J���:�YѪ��m���B޼8g/��!��6m��D;�WJ_p����:�W�@|�<G���g�Zϟ)GJ﬒��ά0I`k���������{����lm�D���b�v���p��.�Y�g1��O;oq�0��?QZ���9�3�{���L&�^�=����t:/���7՚��Κǖ�I��绬����ŉ�������E�}��@��F��HP��}���}a%�{�Fs�u7��1$���V��LL�r�z5>4^X�nAWà����F�3ۡ�%�\�f^��mv=w�KJ"Ag��B!b��
S-7V���v�N8�H���ף��3�@�Y#B ��x����j�-����۹]Z��U㝶�"],ݡ���Ա;��� �@o��%�w���B W��`ڮ�=WEYP�P���a����(q'��@��Ύ�ó��{���K���O�G��am��J���:{�VM�E�g-u�n�9�[Ϯ�V��N[/��s9�a����X��V�P��Z�0�M%#��U�:�ɥ����G -�P�	�lg�&�Q4~�o<��U������P�����6���d�WY<l��*��EFpIK7�%�$T�"-�̢����Z�q����bF{D06W��Y^n���_�� ��B�"�j��SV%�d����ę;?X��U�V���\��T����T@çӐpw�c������B�V�ft^�u^�UxcT�V8���S�C>0T�u�O��tk���o5�U��}R���9n'�,X�'��*���l��t���ם��.�G�f�l��'׃��G`�I���:v�Mc-qj7�ɻ:���BXo��'6������J�Mu��ۮ,���5�Q����1j\~�Sh�t���-�k�Zp���G])s�L��E!�����{!Y\�[;�����%�_=�M�p�������[xwj`�Z����0�������}�:�K���xj:�tuQw\Ra������w#�z\�>����rS��H��&o��@akGG�M�+?c:ta�Q�*�VS��4��}���=7=�d�@@B�����9}���K(���7���B_�b�GxGn�BՉ�\W^ |�N��+mjI��
h��"/�:wupݖ�{
3%o�sr�[sU3/D��G��f�C/~�=΂[�`���/�4�_Pt<� h�]khG��#�(5
�B�]�u��0�\�f��^���u���5���`�h^�ur���%��mR]�/D3�]���	Ny��WALS*������_=�˂���;	(�&�H�	 �M��z�3���_'k^�td�.�-���I<D �a9�a�ζtN7ov{���C�J�F_�O{�>�C4閣��P�p*�>����z���J�^o��5"���T;1-�u���z��vXQ~�`̓웷�m������W�R�P`����D��n�g!���2���m����!�ͭ�����"�j8Dom)��)��%:�폷�əQ�G2���yp����������f|����`���d(�-��6Zm�]�V�f�5	��ef�:��K-Rq^�̨�:v��̃?�g�$z��A���q�OФP��i�_�;�&�.���%���
��*�qѪ�>��d���&Ce��L�����ǨV����)���U2�)z����oM��(���1������,�8v$��D�WUd���̮_���$
�@� b�ʡ�?�B@ m|����~m�>%Et]E��Pk(��r�i�b��uh���
���;�8D�}&(� ��J?�)~���~_��Pڥ���_�\,0?��7�:�x��o��E`���A���MT�YĚ���&���N"����D�\�`/��yvz���9���o+򸛊D����3^����ƞ���bq�z��5<fz�L�Y��*�7-�2;υv9�����A~�:{��Q`=��݅;T%ӱZW;�ᥠ�VЛ� 9ZD�,s��?Ġi~��sC�B����\*�d�l-��W��Dorڬ7
�+��+��7��֯�&���x�UY��{'ʨ"仄�r��˚�'����"3�⡠��[�ꬆl��t�O?�;�S�*z�G⁼��> ��Xc��]���F����'�_B����߶;�DTT����d��Ddv��q��co������a�<Q���۴��	ǅl����T
�o�^�k�;N?��w��5jb��&4��*'o+��[u�K|M��Ё���'�]CzG��K����c����%�&g������&��;�� �n�����hRayK�������=C�X����W�a���KV��gF4>�����۰'���bz J����"��&oN�j`���!�kU����wWA�#�H�)&I��o���mmٺjĆ���K��K�L�M6�=@�J��z
:�0�]q;�s��:QR������^���?���A�Cf��yHx��]�Z����Am�pg��J�U4ua��o/���|6�%�����K���}���\ A��X�F���E��[{��	�&wf�o�2�S=0�yE_h�oXx<�<��Fn�Z���1��#qo�-N�����8v�C�iF뼘m����E�g��6�4�AIBN/A�Bw�g*�l�`�����ݶ�k�@ID��&M��5h�Nb�k�'�!WQ�p�c:���S�w���T���E|b�J}<
�>G��~��t���G&� ܼU Li~pxmrN�;�`���8���cFn��m_<I�k�k��mOJU	7����`��1/� ���ˆ�ET��w�x!xӤ���ó2��6\#�}X���5��/6�ʤ�������N����,��T�bn"[�L��f��~�m:��W�p�I�PT{?:-������ ��]"C�H���[*�V�F·����U3�+C�q?�Y�^����y���j�{:ʞ��[G��>��%#��`�X�����|m��&H�HL�/ߢ=�,^%�np�f�C�NOQ�t:#1@y\eo:��6(����H%V辖?~MH�v��
Q�fnɊ���xPL�_����P�J1i����'a�rW)���<��",����/H�������Dn ����|j"0;J�zN	��%�@k���)R��y�&���CGni%�l�����&�蹾��۫�:�]F¡sꁐ�]�6��5����`�/�K�\:?���p�> }[�'��R)?�
�\泰
2ou�����B�l�W:��b�U�c3���h���1\\S�N��1�^a���~؎��ؽ}�Rq^#���,R�A�Ӝwϖ6�;��!�Rp�����H/�\�f��,P�<�4n5��� ?�7�ǮtAw]����1�j�)��tzh�4t��F��`rfM�)����������[Y���<����췕؇�mkF0�O�s._�7Q}�A���c����\�f-3�
m[�nn�_U|D9�	�(Wz�0_ z�N2�:��ؕ�΂��X�=2y� 1~1��Tj�3U�>u>4��7am ��6(�B��>��O�&N-������>t�P��QM�a(Ѱ��8qC�+�<8���h�eli@S��O4A+&����|໠����f�*>o��S�$#A�<$���)~��s3I�f�ږS�H�^���c�#��Lh9�r��6����0�P�]�8Ӄ#�ax*���)gǝ�g7���R$�?(tn� �P�!�w�T�PJ��]���6i����.���������τLM��U�ܑKvk����K���s��#�:�>8�j�v/}�S,�ϗ�H�B�Ø��@�^K���y���7�v�zO�$��):#�����ywV��d�\�9���y�/ӵ!�sbDU� ����S��A�����ӗ+�{������GH�6��ӭ��W$RLg����5'�>�$+��r��r4v+'��٦�U�!lD �Zu���}'��7�7�ٖw�;ee���cF_H� #Y�"�0�\���)=Ⱥɸ�6�RR�m]�A+�#��E�O�0^^jn��I�]���_ĭ��ʄ7�"З@��>m��f!��R{m�t��w��Y�N���'����a��,�(�ǫ��g�4���-�s\p�u�GҲt�i�4ҷ׺}{����U��TsV��[]J(�S�aN�@�q��J�}w����E���U�~�/�(��n��˼�L�a�DRw�p��������C���΂���KMi.k��m��>�
��eOW.o�㾘�E~r#�@{�D�v��=���Q�$L�+��1lS$����83�!�}��6ƌAP�L�B+/�T����3+(�S��:������-?�/�<o{����w�z6	^����DRg��c�s^�D�r�Bn_��c�� =��[4���qN�ob��%��noG�-�/�@�Q�;,�9�
��)�תb6G~�H�D��NH��Ylm|�%#�%�n�o��%�����r:�^�j=pߓ�΂�W�$�BJO�)>!����G��wV�����MЬ%m
h2F��s����=F|�vrw���vݴ�i]2j^��[e��|�k��'j����� �)��2ԝ�M]�)"px$(*D{�Xx3�����|��|@�`�����d�٩z��3�Λ�M�����O����n���׽xIU�?�z�������ȩS�r=�����N&���"�=_=�t����+&�a2����?_��D!����x6w�ծ��0�{���;v�0��'�CY�fϮ���ջ�\�͜��x��<�j��p�L^yf�������i�*>'s���xY��l��%����^q������*(���F���X'zO<�~�r���|�F+�~��.xMg�f�0�0n�iq�?D�����M+ڣ5}#��#꒙�+�R�Ě�}��ϴ�1���'�:��	2�j&�]�;<Qt�S�k79͙H�~�}aey�a�.����ԫ	���D?o�"?��cV��x9nO�����1pn�ؽ�<��*[���������[����n��{Gg�F�*�:!�Gw���C9���s�N�>_���h�K�k����ѓ���&�w��|(y�P�C^A~;d��	@D��搢p�}��Fd4�G��-�����d�+d��[�&��{z8��W�/��gJ̼H06=�v�,{=��}�~G�#��>�X��DƸ}�,>�\�d�>���M.R��'���߈��Q�(E��èoxIݧ�*0L���dҴ�_��It�u|�V�,�g��::���tW>��e�O��^ 3c�Gr��&A���{=���*���g��C .sؕN����kP�K�MK{v�/�*4Iz�a����<He��b����y���l`&}�w�![4<�"^O�ODa`�{�3C���ny�@%��[�>�����C8u�4n�u.�/��p�u�w�1y�݄K:��ܓ��"��C�um�a�b�� �]A��� ���,��D^�3�@u���ޔ=2;��ܟIC�0{�M�Nu���s=��k�g��~t��|��F�^ty�O<��/�ۯ�z�x�Lf^�M���wm��S�E��5po�Ǩ���]̵W쎌��7
Pҳ|`𚂂�^ubN��D(�9���ͼW��ϯ�~|}v���`��܇z���0���dcP١���
�,4�L��>o�u�ac_�sz�_�]^s���:����υ�L�E�#`�'�J�cz{cSԑ�sӟm���0��ד��Y��{��x�r�^�H7�o� �}翗l5����(�����4�*s_d��}{{�d��E��E�N��x�9� ��Px/���A��t�q˲)q*�8�WY��n��q����y��;��̜̾9Ň�E�p?��g��ㅕo���#����{��ͥ��-� �X!��k������i��<?��6��B�ŷ!`���g�r��*'p��a��:@�&�;j���r{�] ���s�=�7�NV��Wp=��
�'��ӊxI���>���,�l���+��u$�p�i���{-c|G�fPPWP�Ox��}Z�P�M5�����Y0�[W��{5��=��Io��	�!�߇�y ���A��N��-=�O\�z�	o����u�o�g�i�x}�Z���+��Y�TO��@��u�6���3fR�|N���w�_�6�y�J�r�S��um��__� ���ٛRy �Xa�����I�l1M���Hj�UW�r��>�>P���PV���;�#iuѧv/�Ds I%}V꛾��H��5+�7���^J���+=�q��~�p�q�MM�W� �8��>�U���-<l�)nP8��}9�!ea��k�e��L@�ۣ�"�%_C@Pa<�#�%)|k���ly�����^��/tN+P�W�@�X��-D�^��S���%���9Z`��t�g~w>��2;���I{��Gb�Ki�E*���|�\5W93��}L���z'<����WZ��V�#����O�+-���oޫ.;��s�.����&{�����K-r��>��8�Ʀ��|jݎ��ϩo��m6�x8�~[��W_j���+"�����������3����(�Q�fN�{S�^��K-V �ޤ���ǔ��0Z�>n�R�3�����A�D���?`{O����A�~o��A!�������)�<w(U+w�?�7QV_��p͚�&���TC�`��2��� �޽p�:^��m�\�3�WXT��>ޭn��i���uh�* pUa��w�@��p�����IY�y�jGg�}��4Ҹl�Ⱦ�r�Z�L��kj
�j���9`�"[#�^�ϑ��5}6|o�}q_ڠ���2HG�|�Qާ'��-U�e�Z�̽}_�_�Tl���g$�/�>�^����%�3��ISضqا`!�;���*�|{�5#����	:�S��#��b���H��/D�_@d�9
�o'���rxϛ������{N��,�3+D[��Q��]	���ꋀ��)�M�o�S��N�����l��dC��nչn������b���[��5¥C�'�ah�nv���	� 7v���,��	�����7���t�����_[ YS��7���q��ޓ��;�w����ѿ�G����;�_>�W�.�}/��Kr�;�w����ѿ�G����>��:d������삥��c��bc�n<���NӐ�&g�pq�KK�Q���K9�<���ڒEG�⶿M�� !�ꧤ�'~r�|a��x����KI��钨ە�ݮt3Gnp�m����^z�7����K���mPT��r�}�d��2t���=v��*{U��Ap�Þ#�����?j�S���ߔ���7�)�M�o�S���ߔ��)_����g�M�G��oj���N��g�t�R�}?阉��;7����uG�׌}���Ds���r^nU�ؖ�`������,�)?��˧��a��|5Q+�ß�{��8�m�����?Du��b8
�c�M
�
j3^��(Upkt�ޞJ�9֋�iz����ogP��ol4��)(�����;�9����:�=��W��g��YyO<ja!6iKi<�e�]V�Ս)i��,sg95�/��������5fސD�ڞY:��(�7���_W_�&�415�k�f[�i��n;�Xx�UG�?M�� 0_ś�fw�7�\57�R�_n���'�%6��E���YOŌ7W��d��3��Db��^ν��j��9>؀�
����f<�X3����%��X��b��g�� "$RL�SH�wTK�Q����?p�|�5����������]M$-t�ǥ�ZHz�_<:����W$����ʝ�%f��ԫ�o�%�jNXwq����k(��qp&j���8{$�a�ps�Th��$Ĺ�H��G��r�Ֆ��iq�{��E[-���'����<Z��f��U�!�a��T?<�8�̜as��)��cǎD�sM%�&���b�����L�V9�;�����$��"�V���>��Q���f��Q��	.($�Oo���͵���؝���,VcM�۸o�o"ی�VX�czg����о7e�ξuُ����f�E�`9���]Gq�>��aN�-FZ��3 ��4��8�Hhc�)['m2:y�%�mT�d��u���q+�	��z�O�S��}qH3r+�ܶ���-�pu}��z�1:�СIm���?��=���j䯙Pg9��^������{�%:�IKTg�e2�F������ԛ�iWu��-a{�m+2-PnWn��	٪X�-ߺ-�S�������1)��n[��[߳�mf���MƎ�>�l۸��r�9W8k�F�?L}�J#i�e�eᰏf�zMb,��P��[�飽�7���둑B&�o^~�L���Z�N��ά��v{��T��k͊�K��&���{i���_N(�����1����z��Kn��1c�y?��\��BYw�%��ޅ`�=���3���*�ө�y��Wfr��g�:T�5�n����fI�|q��r_6�_�ܡu�`�i���Q�[\����/��J�@{�,1�57�Tm���R�w�C�.�
++��<ΰ�\y=��.�Ƙ_��r�ڊE�{7�կ|�����A+��"0���+!�:��Io"���)��h���b�3�	K�(zS>\<��
���ŝ��|�嵡�����3}ȥm�LVRl+8˝�Ě�(g1���Zל�%vC��w��W�;����7j�c����8����k;���>�M	��iV���#Q�St��ҕ�#o����q�q 0S�ɦ�o��A����=c��@��;���ݽb���
���O�=b���+c:��iV'F�(n\ǧ�%�/����q�<o(�C����U'�MƎ��[T&b�EU?�عf3kt�t��d��j���Ғo��ƌ@��H�r���sGc��e̓�+5h%[q�?��i�G�ګ��ҫ��3|UUx�R[^���,ǵ���:̾>#�RWR�f���'CzG6$������l�\ΆN��G�M�úu"�������JW#��5�ւcǅ�'��j����c�6�����7���O��dJ�-�{
yAH���������?ԽwTSi>ꌟ�,���f�(Uz��.���;F$t��"5
қ�;�K���Бމ&t!� !�s�03���u����Z�i�y�w�g?�>���`������Xxt����=�eР�SO�d�'K�"��o��<5kk+�ß��4�`���Մ��	�ZVah������(������a� ��m�tNx�f���+�Y2��Ӕ#,^�������V�j=��-D�$R
��Ï^G'PL��� ��ǵ�Ҵ���(���'L��������ܤL�'ac�u�"{zz����	�Q�Ͱ4���^��, �!�\�8�t�qN��|�XQBG��/���z�������璐r�+{#�Q����F6ܧ�� 6��i_��%�����ĕ���>�f c�O����X�pR;�އ=�
�?��,�h���v����L�,��~d��D�>���"�#�U-���s�[{追�~�\~�U�����y���^2�20/��%cK�Q���m�|����W��_�I��f*�B-%�]�c�~|WVV�K�W.G�R<K/�c8Q
���ܝ2����Q Y�&���-�F��ԏ8oC�
�.��^j��04qWG�7�s~ Lݽ�C[Q|�������xzTw���Ķ_�߶ �!���!�4���A�7�����s�ec�����w��'0=i�t�{��R�|�[�q~k�������+���U����:C�Y��/ɴ��@K=��w�hU��F��BXZ�57�X�aЉ��CIU� T� "<���u���PIz�l��RR"|���P���7��#�N륿 B�]�'M��o�7tg���������Tm xV��v��7�j/&{��'i�I�p7az�(��P��!��E�^e'�N �r0-�X�G1�\j�}�}�d�))2A�V�xq��.�����*�A|9�"�O��&{�W�笝�-ur5۫5��O}��s����B3�P�0T=nڸ���� ˽�jd��b�4���"�@~u1�.����D��UTUz���W���B"ha�U�̦�yu�ӹ�͓c9�2zCd�ԖR�K�ʟ�a����e06�w&�G�(kw���EW�� wb�/k�S7Kqk���������8����,�1�����ϠQ��$��o��4{��o��/�=��=xŔ�sU���r����¼*�6"t-��4��tTo9���!�Q�,B��o�Iڣw���u���N�7<g�g�;� �Y~X�x�H�?��(�/�˸	�4D�'�i���h0#�	��*��<�JQ�zoٵ��Q����;lܮ�RA���g�8ҍ;(rE%e೨�c��}�G����&�(wj#��m���A���w��͒����dUG+�s�8�$Mj����+q��wܧt�	V��M�I��lh��R,��K%�Ļ�ڀ�E��W��{�d�Ǿ�]"J���5����0P�V.n�eal��Q]ߵw�Ta��DǴ���3(�ٰ&�%e��u��^U\8����2��IR���Q<4��X����3O>K���I%Wl�1���[8ք��8�k�w�I���w#o�
�^���9L�<�_��������߾�'���B��C7�E�逥��"���{}���6�K=��kr�)��K�;%�Τ����z�� ז�-��}3&.�~;͏'f ,�C6/"�>x�����:��?zd���e�o3M)]�������ҙ��Qޘjt�Nl��`̰(�;+K?0���M_�O�B?4g�������W���0����p�a��`D8��/�jĂC��;����J�n�n��kHr��xۂ_���yb���c�]K7BBc��9RA���]�G���#Ӹ���D5��v�r�\�g�c��?��sL�V��� ��3�4!�pr��-�p�0b}}��A4��2�~��&�<�@Ȭ��x��HVȠ=#H�3���]��χ "5�L�R6���nx30�O�F��n�s�$��#\X�˗��e�x$�!S�E*�bݷШZ�J;8��~$����f���t���HZ�󁦌�t�/��?�:l��Ô4�#ۮ4�r�{I�uvu��1��[IFM�Y��ye��M7��?ى�汹v�>>x�<��f%�Ó�c��d�)u�NI�TFA|�z�J���C߅{��E��4(�+���Ijj��<3B5�aqDپ�๮�o����@����l��&7JC�S��5[y
��@?Ű��Ej���3|;*��齜g�Uee5�cR�r��V�9{P����Q)O����,��;KZ2��B '�Am���&n��gi%�idX�B=3��s���j���x���{B�{B#L��bU�Yx�<w���=U�^��D���N�����M���-䖬0�<5�Np���!}��T{)�-S`-�c�g!���9�;��4������K�x�@^2e��?>���}��R�８b�4@̈�k�8W6Z0�,�eS^��V�_�����N5�oajޗߋf7X�	�n��/���(*#a%�}5A����\��OW���B��FMF(n�x�����?B"'��~�b��cb����Q��I�r� 8$?'|�*����I/�@k?�µ�Фg������D@�ls>�y��`z��b�>>��}:�M�j��b�oS�����41���]�����o��Kb�Cf�+I������z�� b�g(Œ��W��}��8C~{9b\\��m���lݲ�{^��s�+��g_"�v.� +��.�\�O!l����%���|U�Pb��匕��3ឦ3c)�㠻��ݼ��|�RC�sU>j��w>����":܏I+>'�XV�6U@pL�zǤ2� �J���ƈ�*T�%L�t��9���+T8��ՙy�ʬ�f�r!6�E�KqӁA�	C[��%j{O�JQX�Y���I�O.��N�Ҋ�yg�����lE��S�#Ñi���LW��:�XMf���D�>F5�����[����ѫA��f�ҥ��T��J��/<�EI��76���ȳX*8���� �e�)��F��9�����A�=��a�aZ���Y�����_�59������_�h�Z�B�up���:&5^�jD�]ܱ�h�~f^�6zo�9f;;���S�*.ư��~�7qQ�е��r.�LF�e�����4��av!6rB�!��_�����>	�?4��iڙ���?���1�����t���6�7l�����%6�O��X�a덾�4��dhU౯ulw��u�4t���&cD�8
��b?B{�����#�	�,��Y�S������"��,�q�w��>J�K�`���b�J-S�J꺫C�Ԡ|C
,��~�?��{�,jx��ᑝi�,�>�?$����#�P(�X� `�\��AU��:B+P�-f���r$W���s�*�[M}�s��2H�L�^
�lZ]~b
���HW/U�`\w���� ��fwt�]9�W|���^�/U0���fOí�����ݔ{�Qb�2k�=w��P�O����[K>��@�Z�Y���Qh�*�r���C��-~�Y$d~}6��W�"q��j�mD�=�`�2�k��\��4.%|N�F�.�Ov�{N􆡬��,�h�8�6{l��R <ɑ����XOR�iz�^O:�B$�dg�7��{��C'<2��T����n�+�7$
����Z�?4@M�qE���1���E�RX�q_İД���s1//Y�gߙ�ߊ��Z��vI��ke��z�1�Q��!U��yKu���ԃ���-|���
��4�ȟ�y��@UNr�j�]��@��&Z~MA�-;�i:�_��K�Þ�3�Q�n���4�f���&n8ױ����4M7�~�MR@�.9����]gqh%�g�̳��݄�rV�?�f�T�M�e8�.�n�N�fg�G�����	l�M�������Y�h����DZͰ0�#g*�an�uB	!U�����r:����aaL�p���t�vaW"�6��_w��~����I�m��$�i��B�K�F1Fl��u�i�>��s^T��/��o�')[��~5������g�)�J���~l��U�V� �GMm<���k`sI���ٕ���*���R[H� �MӮ�tJ�Muiy����[��'����m\���<s��lI����6�;R��<��n^��>�-�4h�5�J�u�� /����~)7����H����n>���2[���|T��$P�ZL-�������4hڍ��moH�dcmg�#^��5�����DuL�~����1T�o�"�3×�l������Dk���FkO�6�7|��/�g� �k����a,s=h$n	���b�ᷙ�\��Y�J3)l�w,-��Db�,���r���=2S��'{Ol'���RA��O��֟�0Μ#A�L>v����3Lqg1�!�;��^N���WSQ�#�!��'
��C���4�!�����(Oj��ᠭ����c�n�࿅��>�o^��!�`�d!�',��4猊�ü��x��9�?Ld G�֐��O�œ{Y"î��wi�M�����=����'(!3��a��)�=��Vk����in���J8(*����l����O��eP�utt� x��+x������{	��pN�l�>��[�+�sD��ՎO�\D��U�{���*cz'����T|�%��pOM����;&�j��e(�˥^��ֹ�43�Oʰ��a�..y� �-�Ǯ=c�k,������pE�H�Kբ/�D��R��z��\Rf<�v��Rg�?5r�Uq��Q��N��|��kJ�J��~5ɝ;Jq��g-=M��s����S���~S���˾oΜ����/�OTkp̷Tӑ�Hl1�Ҿ8��{��A��Җm��)���♣�)?1�gg�x�L���ٝq�����$���/��@��|pJ�Y�O�f����gs����T�m�Ǽ�E^W:�ʅܵ�-Q�l��rUU.Nnlt�/ZZ�9T>����k�!�v'�$\Y���[�����Ɓ�׺wVuP��ʅ��7�N࿡�m|��h�4��d��U ���[�B��8�9���<�U�z�������6t҅̐�����ʦ�M)��}��Ȼ���X��
W�]	�k��
��/�8i�2�I#�6�%~�u�8Z�I�x��NF�[��7xS�ZHp�=��ɑQ�r!gh�i9�6�+Cf�O��/��E0s� ��g'l��/�C���"�sQ5��CaDYv<h�G~���W�y��P�Z ɪ�x�oF���8�E�@N��c��������oS��	�[��?K��� ��ه�Ug�=_ީ{|0�2s���uڎa_I�ll��b�gU�-��n���I0h��gާ�`��o�%�-��q��;
�I�����8�����_~�?�¤��Va��X����"	�7����'��n�a.�IP�A�9��#ʲ1��j�O���>��� O�T��Y�G��Lz�O�A���B�����՟��w�E�L��"Ot��_��5"p��?��Ν����N�s��٫�%H}��xA��&h���|��������k���G=�!��6i5GGwD���:�f�@	�%����"]P����|r��wk��B�l�G�3Y���Щ�>������}��v@��/`w��b�k9�����v[������^`r��!ەvGC�w'9O�pw��ʄ�E�jh�_r+}
t�L��vW�]�v3�Ѧ{���-_��}�_/֨���U8?�-��:�C`�Q�Wi��A����O�m��Z/W�
���Y�{�9�����q5�9�����6�0���ߓp���Gc�r�C�r�r�� �m5��C)Ϟ�ɋ��O�kf>�`ZP�W,�����ot�!9s�J,��@@�u�D��-�8�ehqI2���i��ncExB�L�j������`"p��'��SkY��	⟂�}��A}~S0Z~E�5Q0��7魩R�8-J6����m<����pYh'?��pu��X�ʡ�F[�ENxN�V�q��o��d���V4�=#��C�{%�@L�S�n��{��H�˻>\��|�}H�W~����0dI��կ�sB�/���4q*�q�3Q���dG����d�"}�ʁN"U���%$ps��6VZ�3�M� �hA`�}W��	��8����o~XFA� c�(Lb�iP�+zF��s��l������\�U��r��1���`�r7�4�.5Q�Hb�9~2��tZ��<���j��'o���Kb͠���(��� 5��(B��U\�L�y�y�+��"�egN�\ H͑9���y	���/dK���唉
��z�{[#9$�Vj������|ʵg~��/j{���Q�>;�H��Ȥ�{{�3B'���.�F0+=7���a96�_1�x����������{���je��N�D�K�r��*���B�o�j�j_�q4Da�?��3�݈�}�VQ |��&�~��T�6����@m�G>�:�>1{ڏ�g�V�8���Ŀ�%��UR�.������\mm��C�B���_cr�Yh�޼qY"U�I�RC�L������l�l�`&����&��7�֑ͣw�rzF��5�:�yܻ�8����lK�yj��VPj�����a�Դͤ���B���$��nG���c^��V���G�}8ea.�\�|v�ˋnǖ��A�LJ�s���llX��J�6y��۹Q��ڛ�)߁�w���tzЧ�澛֫�"&~��e/_|�m������JUQ��;\0Fڍč�V,�`��Rv� ߂}����������Ȱ��t��<k+����Sa{P��o��tHF�{�7!�I1���@��뉿dI��:3�c�(�հn�b�>P3��?P� ��g8���~g�����sb���	r�r�(Q<D���NUL����3��i�����4
��'�f���=F��ZlI�+�5��^g��,@�DQ�U��W�ߩ��>R��7w�N{�FT�?����<K�9*����"w�i�$����Z�%.�ފ�9\�)%0<5���1m0��m�bz���.�6'��hz�y����vc�t5�?�]MP��.Eq@����q�^l��s��MX�+���s�	Lˠ$�����/^f�����$
��2uW^��B�u�Ʒ���`���o���.�Qz֚���R��fx_�w��D@p3�9<6�c�P��ۣE��^�Å�M��5�.���Lн�TQ1� wG'V�W��D��nEt�6*�9��"�D�ˈz|�Q��\ڮ<�-����`���K�R�d`؁M���ؗc��&³�2)T�~���\�:F�1_S�t��4����1��l���*E��K(?X�����P�Ǹ�<(�W�<�&����- ��;�����	��+�9�0��7�/��W�E��J�̀]�d'���E�m�	2�� iNCw��c_�X��ŝ�R�(��*�1{�"�����\̋x�񅊔�0�6������>99�^����DAU.�0�NC��PQ�[����,����eZ�vƳ�3����W�o���Q�IήAV��D\�G�`QZ��½Ә��!����v}��H�wܾ7�e�� A�?�Hƛ7�]�#xW}��m5���鿓k��7�:�ucR�j
,��)��)O%���F��m�#�����~>��p�k��S&����W�&�{F������yv5�����<��J�/:��4
�w����@\9���~Nʕ�j��&4,�e� ��a�Y��0XgK������]��j�L�OX��QA���	�՘��[��LO�v�Q#�<}��  <���o��Ȑ��ߝdF��$���{VK�K>]�d��N���i����]~D*�bd$�'do+��#h�G��uH��d��1u�DV��OR؝ $x�|�`[g�ɟ��#�=�G9��X�������W��fQ�\����m=��`���S�(�[�^�)\v۠�<Z��ﵞk��50gpkD ������Z6�9�b��_��>�P ��-���	�?բ�$5�P�`wn �c�{����ވ���PGɷ��`d��޿W���v��fR��]w$�e�5 *�;z1ib@9 Ȁ�j$î�OT�i� O��ۋ�i�O�A��=�����i<2}�s�X-�)n�K�vr���С�U���A6ﳅMT吉�I�߫;�un�A��N:}�׏?0����݉��܀��c��F�QS�$Bˉu�m�*�~�V�͛��k�ar��F��z��=HRV��-���ݨ��[�t ��Ul��~9ѝ4!�W��MMA\S�҈�65�ڏp��`	$K_� �הq�G�F!��܅�lO'V�M7 IeO��XI1�Su� �A#|��;�A$�ߊ�o+���D�z��T�L쥬3��xd�tc���ّ�թ@�;���ܬЧ@]3��ؘH����IL3�P��Ȯɽ��(,��]����:�2)�%�����(��@nM\�d�,������@FK.�'�Q���|q���t���߃;�M^����%��w|� ���cS�`�c�b���gw�(�EWͥ[��:##8
��
�)TH
45;l+l�+��جW�zK��nH|lT�6�i�K��z�Ϧ��gT��~��M�b����}���Ԫ[U�~�;ao�ԋ5�k~ �L���1��ՃG�HL��� �I>Q;��ҕT������[�q�E��� �aKM+�w�\&���v��Q8�I`J��k��.붦&/��]��BYw�9ρ�3j�*��	�xޒO�4��k�7���]|d`��Z��7��`�I�z��I���T��RsI�N�^wttZ�Yk!��o�Ǒ��ҭ��G 7Rn��_	J��r)!�Vh;�0���~���u��O/!��]﫩�7�)��!�M�W��d(�j[�ITR����k������V	��0�֌�i�z�Z=@�Wı�x���?��Ş�W��_��>� ��AW�Cczk��Q �Y���fa5�<��bF�m�+�j6�Tg�p� =�w'L�}%z���d:�Ɋ�Ż�C����0B�s7�_I����{���5�.k�&�sg������$p:�tc�Y�-���֓����I�����|$[{�7���� �v�������g�`�	a�r����˧�w���G\4��0��S�
�~�J6w��[��	tZ��
�T���0O���~	�<O�3\�~{Q���	d\ �V��f
��
���CZ[(�?O�OTT�fˮ�b��0�E��"�긊S��;� X�R<�$n
f%��Y-�M��(u�ӓ֫�>�{��a�R��F_g<��e{l)ҙÿ �g��qO*�=\GR�8K���"Hg��gK�]0BnM�"��Sju
 a��6x��l��P��98��������i�=�6����:���
f	���\���,�n
u�R�4=@o�H7���|��9�_d���'Jn�'��dp�V�)�͓����j6��k!;���'u�.k��#�2}��:���Bn�h�ܐ�'^��`�xgM5	����Z���Ύ�~'2��H�<��AK��BO�j���t�Q�	C�5���pb}����t#�]L��ÓYg��_�)�����x�C,���G������"��A/��I������� 	�#��VI��)hM��J�	�p��)�a޲��-|�<|�
�Kr���~���5�	1�][(m������C Ɉ�?��'��" ��$;�縬^���=�K��@W�$�R�\ٽ�n�^�J�kw3���`Z[g�A3�6m��&��´Hd�ϣ�,μӕJco��Q�pQ"3�O:�	��@xUgG'f��$؄��9��!��O^ f��o.2F�=P�H�/���.Hټm�~G.8�)3��S��ጴ`��߀��>���7�9�\�>U�no��g�(������w��G��E���S�ɭ��ߋ�b&���X��@�#Ψ�%N�V;�Ǜ�@��d�,j�Q�>&+ 5�N�}h�����F�'i�����+���=&Q̉������u�EP�z�*ɕR�9��$�3`'� đ8�V���6���n�@�4����St�p��>jG~�86�ी:�0��)jGKu��7=,��˩D�bfzN'�U�I�s��v吝)H��ү��(t�9���� n,dױ�8���P������0Eズ�5�*��dH�PN8��VS�\�fWbZ�L>����)�8�-���[񰂷4����(h�G7��b��3`Y��z)�iP�ӓY �bI;���O�W��1�˯a�y7<5@���8Z�� 	R4�����k�������Ik��=�|�0^��gu��V^���,,�]1��^XԷ�CnVvf:��]p����~�����`oNठ����)P��NST`��~�MPw1v������ܒ�7ݍ��\�S�s_J�-BhE����̓�����4,Zcg���5|�^5�),�����J�M�"(Ū�NS�*�A��+�pb�i�f���������4����	S��^ �5&Z�,75S�W��ɗ�4|[t�� *��C��`��z�3�W�
\��w�tʕB:��%�n��]�,�J �b����l�.yęDfk@��e���Я��u��������j&�H�+a�@�����D�=W�@t��e� �IQǙI!��	�?p͋H6�7gv���ȒЖ��J��ϯ,�U��Z^������ 
����Z%���X���>)��*r H�������i���U։��(m���Mw-�Np�g#��՛���͐�rc���s;�Wˎ�f2�G9�;ϧ�O�&�`�;�1�j�h�S�oSk�J$������m,@t��l2��2~��
&\��	����c3����4p�����Z�� =�OrŲ^�vV����3V� P����0�eP0ͽ�St��U`����ă` gF}�4���i�	٢�Y�"���x�D����q��ĭu�$fG�<�CF�c��)�<0�O]x`�$�Vr�.�j����N�������I�����z��(C�Zj�+#k�#����_���� �Pz5kh�3�������9��X8�,�zFb��_��s�^�lԙ��(@:_wwUsG(pM�<{%X黪���W��r=�7{< �����#��k�k&R�x=5pvk�ߵ=���4jZ�7x��v���D�[��qOз�d�L�)�G>hx�J�e��	�✀���(.9�sբ^E���E�:8�����BB��h���n�Dv�I������S����l~�'��O�͞L	풔������`}�϶����~4�l��	�����ȽnS�Ep9����~iG���bgȕnHB�Gf�V� x;��m��h�p���,N�H��U��p�|F�ĭ�7[^x��p�w�	�}@�� ���ހ��P�ۊ��9d1nR�-O�pb����;x=qށ�/�GO5H������p-�tHТ�~�d�}=!�_��-K��H�=Mޟ�N���5�����>�N}�|gP�'A�"��b·/S*���ӧ �#HA�(�c�
���L���U��R���.)��m��m.quل�m�I���zt��1K�)�c�N��4��k�⿞��Q�z��c�H����2��yX�j�Hχ�=���̤a;�X�uY!O3(��e1N���3�$*-=��W��]J�# �1�����W�ε�XiT��t���2Wt�2�FD�*�e5����F����@��v�KC�+A�ļ����/��*�D�c� ��]P��u��������&+!�����:9��s1 M	�J8��H�[�����������1[��a�۫l@M��%�񙲍P��6q�k�+��C��M��YBMY�9�jM��Cs��,�fDR�u�e��>�[�V����it���ePE���6��^X_߱���V.��@����҇�V��S x�&tC�F�����aZ�8���T���]�nc���Xd��r˻��������U�4���`&��)W0���/��T�T;�^s�����3�A���#�R�l)�bp��|��Q���	ݘ�� �T�)K���<]�vg��H��o[��k����
���X�%y�G��W1�y��3E���"�әpo9V��og2(4f>x������ǫ6���O]>R�5e�K{ff�tN�L�t�iwimv����^���=�'�6W��&'+�D�-;뢢��
�:��	���y3ߪ9�R�d��d��Y^�H)��������瀋u��â��Eƈ����ϙ�[��5RN���p?
L+\�nx��'���R�ߒ7ݳ]�xx�P��(����~��1�8�2�v��m�&��/�H�D�J�N�]P�d1�0�-1��k�P�a�=��Ҡ����BX���u�$3.Ss� ��b����Τ�فI�I�1���
��Ơw�N�㰷���r��T$+�@��y�w7W�5s�\�Q0/}ƩR��Ƚ����)͈�[K\�ƖeBnA���$6i/�?ϰ��).�u�L�rj8�p�죡H�o�a����������'T�*-�hV+�I5(�"S��B#�'Ĵ~"��J��q��m�o1�!TJ�x���t?b��6�h��-���\����K��S�9zuz����jbEFE���3���Y�4K6�������3K�1�2�̴RwP1�-��P� �{�����������T^-t���$�Y�Gv�R�d�y��e�Ԋ둖�e��ZpM NS�9�T�8s�r�Մ�a�9f�W���+S[e��ۘ���"U`i�b�\J�Xz�[�;߽�7���6�{�#��a��j�Uz17���O�z�5���>� iĨ�1��p2ݥɊ�D%��J8~�����)��.�����
b�U�_@���c��-������.,���� �F�~.�|���~6�$9�M�|�>��]��a��~���4�6�ߍ�lS|@	�y^ON"@���(��=���o��WhRMbrm@KCl�0���SҎ>�Ft;�r׋��y���P�>�}2�x~���!��|	����OmkT�O�&_�g�c�:;���)��O��h=\N�ÿG�O�V�n��ݰZ
���l�Z��8��(5X�8��,�E���C�bK�%=��HK�Jk��Wxo
]C��A/h���bz�h����b��*�/ۡ4Ե��r9�٠�Tt1����Q����N�Ɖ`��^�rMz��<r�b[b�Z-�ns�E�Q��O�����#�=�1�+b���"񚠠 �{ �VM9�J���"��Яw/��̄�j!p�W_��c_$Æ�Ћ2���n�R⪪jG;�8����{��W���#�{��娑@��?�;�~ LUE'{m��̓��	�`�+��hѻ^qd<���0�
h�v_��Z��Ҝ�b����$72��}H[K��'��;{}"�K��M[��S��=��9�{S��(dJ�6Ub���*6��e���J��[!
�<n�b��.�Kw\ƾܛ�޾ݷL�H����f��s1pi�&p4ר�-�?61����z�7���6.��e��>��r.D�?c��d����@�I�w�0"�-,�5RY){)�����_��)��a�b�ݷ�Y��m�w�29
` (�F��4��ȿ�8��p�eha�)9���X=`�̵x�Ba��, ���FI'�m4���Jr^�i
����n�j�]k�F8�ۦ��mh�����zr��s��50�31���Fz��t�����L�Ϩ�>�C�
s#ai�f���us��yo�G]z�͊�JJB��e/{n��*�}H.�n���H���v6%k1��t�X�9����-����Ø8(i���@};��������P
���N�Q3,\� 6�N.�O���4�ݽ1�����m��hGBx�,�@��4|[u|0��'�S�?e���Oef_�-|ҒX��>8JO DmX��PN��ޚ�,k�녜5+Q�3��-*
������`Mw�q����D��	V�̓'\n��̠;���-32p�jq�7��(���1ȉ�#-�'\�8���g���~���A2Ƨ����j�*}5&e�!�P=�C��������̝���fϦ-K����|y�V�,���GNv.����Xٓ�5�����ҽ���H�@6�(�Ra��]syugW�LJ���L�ƦШ���9t*�9��b)��В2�TOm��~����z7���z���A�5�J��^I��M�><���ԓ�p��;-���(�ۈ,��4�42�U;]�q-�����X��s�ʄ�{|�˹�"��v/UP�K�e��=�Ѝ�\��E�}���x�k�t�Ec��U~�t�����彘���Zf P*N�� �&�\�!(R���	��Ef��=;�����Y�ߒ�-��ۓm�x_�'�[m�0��1�:��h��@�z���6���|���r����RI\�N w3T��@�~Z���l����!.�O�}�v��E����%�� w��P�����y1����;0yƂ�"��(�C���8�7?��k"7ҵ|���KP
��#����4�QV�sv5 �	�b�pҶ�����k11qH5\�_�*�:�
ױ��Uq����G��)Ե �� 0n�܌F�6gr�]�r[���IbE������U��itsZfw�l��<F�7��ঀ�A��I(/�r�����Yrv�����(����7����4V����P �n* �$ ft�-Ѹ���<�NâeK�_����$6��䵓;P�ê�M�K`ث ��T��C��םp/::�/�������NBJ�%r_�	X0�(�ŕ&�j�fhXh��� ���c\շ9��Fr#D���}_,�2����n�Ի>����.���d�� ('�����7Àp+80�W�5:i�K�ʝ�_t��~=Hc��p��>o}�!#��Z�, Jl��� G�ܓ#o���1�Xס�'�Øp�����s�QU��c�$��i���?72�o��8���2���Y�:4����`�Uˈ���������1A��԰-�x�w�f���e�X_����)S��$�-�ؾ?yO䒅�ôP��Y�'�J^ѻ"` �(�/﷌ơޭ��f��Z�,U
�vT���[^��0u'�j������JS�F������9_��tϮ��\tټ@Ѽҋ�M�IB�ˮ�d��%�K�2�R����iur��p�+�������A]��)��+�[p7&�}�;��X31��B�i�w�� r�5�d^w�n�)�G��&a�����9�G����[�d�(i#�u$���/�p?�\�yiϭ4%��*�Q��F6Χ���󣏢]�CtT"����ӵ�66�� "���e��rv�t�;pƌ�x{��Uz$Y��s,�a]S�d¼Th����?5&����
z�3��� �T�?�� ��@��#nJ|-�#E��s��i��N�)��Ĳ��U��`	-��-ւD9`��Aт�wB�6];���R�����,:��!��kn��R[
������?qauYU5�&�E�!��+݉�&=�I㍷�;V]����;�}�iǚ/2�o8�n��� �-���z����=�Jeuk��ZT��s�F�m����/F�P�Hk�qA�� e���W9�^3��7R5o�$A��ʙ����v�b�*��0�}6��}��6/l?\?���l�᎝����A�ɳ��n0e7�7\V�m�z�E �y��t�J�$ٹ����\���`�"�}Q���[�~����p�:ⴟ9+��4������o�,� �ftP�1�g���n�Y�?�9[�j����r�z)B��h�F�pYM�U�����9So#	�����Z!�^�q�-h2|��eN8�|�c.���?�=Hìu��R�	�������%+z=!��V�����SY��لNϸf@�r-�Pq�}w X#��"/-�§��H����^�,EO����3�\;�,�l�[�a=liD��d���!���zjo��B������т���՜�=bg	:y�B)��-F�*��}U!,8xM�c@�G6�Ƀ�w�?;�V0�S��ʪ{�W���>s��R�����!�y6)��%$E�� �ߊ���(Ra%��n�Wv�B���yz\׮h�;%���l� PT=�L*Er#���pI7&�#�wӬN��	���� q�K�NPO]w�X$���Nl�.�|���z5k@S�7�0����eN�x��M@��䬱M��Stog�N���}���kO:g��^`�F�D�&��˂Ǐ�o-���J��C��#vA3D�;�W ��lP��t�`l�&�ߗ��x�n�$���0��G�G8aPE� ��	�P�R2��a��݈�|5-�o�PV�?�jYl�"�gb�sLI�4/G���Iu7l�lM�ڃ�z�d��/�g�Ŝ1��20�yz0]=r��A�b��~u ��� 6���бF��Cr�R�]t��NF��~K����˥��1��Р/+�m��7�!j#}���#����Q�4H�>�+(]�d.�A�+�,
 6�t��m@z��S#��5�L{��Ƚ�+w5	��~�Oa=r��X�	mҷ�K�����5��BB	@�%�g_�-i�w�2 >�[�nC7��\�qi��&_[c?!�/A�~�4[��������]�8"o�D�Ec>��ӠV�񇞿�n?���-6O�>�=
�{ǡi,��-����� ��=S���1B�!��ǆd�NM���WGB]�֔�ҋ�K���df8)��h���iPj���'q�x�m���o��R��?�V�48� ���)�>�Oӓq�~PN��<�2[��Y?��də�erKJ!ś(�,}��q��g�72;�9��<g{�Q��9M��+�ө��t�W�i�V�s��AIܨ�\����N�emX�tɯ�k�����Jn]P�����I"OC���g�u�O�ۛ��\:����PL9M��ʅ���>�{���Ț�z���X�{=c@���n��5b�\�	���&��M��ؖ:J�R�Y�.�b(�4���Q���"&|����~ʿ���8�))��,�P��9@�%�C~��[{&\i�%�mW�	�%z��y�^+�:�P�b�PP{��~��k��Ж�(3ZOVڠm 6E��ƶ0Mn{�ߐ�U�*�q'�P�b~6@a^��Jo��C-}����w�e�6��-Ux{�y����l��M8���������#�<s�,RT`%g�V�/�3����~��V>v��8�gP�(B�т��A�$������tZ�U�<\������p���bw�`��iX����� d
�bƷ���Iw�J�����<i�a�F{)�ݻQ��9�#"�@KF�U#��uꞩz<�b�0� X�~��C�Ld�P�X��4XĜ��n��a���M�t�)ֵ��LFX�4[
��A�Cm@q�����S�VP�#=�[2��3{T�!�����kroy�WN��I-�'��A�����N���J�����-�%�s���!��4�ŹY|��:n�L6���?��^��HM�&!c���R�V������LM͓QK+��.e����>VKn����Dw��'���Y2��A��Gbz�*ҿ��)��Cl��3���Ra����u���P�HX����e�@�}�;l?~JR����텈X�!�	��c�<�={���)�/�3*�d[�E�qP�A$IV�MlP�YB%(��$�d� ���@rlr� ��᫷	:s��q�����̑�ߪ����޵�:I�&���U��K�]#S�ڲ�v&�^�W�[�W�ڛ��@b-����o`-:���R��^51��G��^l��F��ŔJ"��S��6L�K4�,5�|�hkgRe���LM�of�Md׿�T�V8a;̹P�+��r���HC9(����VV�Ȫ;� tb�P}����@6"ⲝ�ۮbU�v�=z�����	��G^��$���(���z�夆_4JVu�uT�I$�mdA��W��>�^�	��<L��r���['��	�)�>:����`uǊ�n�BF��N�S-!06�Vm嶐�.�V��yy^i|;��lS ���-j��Ĕ�cY��]
ȣC�����o��7�l�D�G^�q/�]U�{�=��(=4��]fC� �C����Ei:I�Ƞˈ�N�ƶBA�r���J�V�U1�:�D�U����(W�e����M�1��I,Sq�|(��_,��c�ҩ��W�꺛@[?7���/fu����T|zI��\c]�O��.�f���Yk���./ۺ{���Y?%��y�:���Z�t���]stqY�rWI���5��[�t�i�-�%��7����0?<�{d1hWW8�V� *����T��Z*�j��,��`���&G]F�+�|�J��ߤ�����F���S�
#��u��5�\[�tm����x�A�^24�ʟ��r�`@�b=�![�6��)����#{��as𝕤���lm�P�hR�����C�O�&`�}��D��W�Y_I��$��L��m]&z�>�1L�f@�ٞ-&�i�	oꏯ\�v���o۝�q�4`�.�t
����P����J=�l��T��N��]�5�.uʦ��@s>���v�
*RԄ�IAg@E2��� D[\q�(�x+�^��p�d�(j���� 4��|�U<�K�F�ToLn�������9c�ی����3ܪ�N��9�	�&�Ft�90`u�a�U��ЯuS[�$�T�p��|\2;  �z���p0�T[�uh�,�t�UƠ{a��s8g�eu�LH"PO6���\��hӶ���6��\T6z���v[o~���Z�\����L�n��]�"@��-6��A����=��!��Ƿ�^հHK�X��!$�!p�{K�s�V��Cݟ=��a=�)�ҽ!O��,�us�4�@��A�;�s#���~S��إ���5�ߏ���5I_���*��JO��]rm���p�|�s�K�g��UmV�B/���#=#p��-�fн3�%�.[����ڢr�rΧ��]��Ռ�`=�MAj�����n�0�����uӕ�v��zغ�ܬ���HA��.xǗ|�(�8�B"*�?���j��	ڧMl�D����PS�?m��CM���m�\.��q߁j8�r�	E��Q�P��j��3�+�[@Y �o(�����ss�h�6�x��0��@���E��H�5���B�r�����W�����3��GG�:��u�ſ��^�61q�9Ά�v6�'�*���Ҥc��B�2��L֎���P�0`Ư%V�T7��Ջ��2iVC���d�kR����#��"�q��izm;W��=xS3�۪S���G��{Vo��_�ze(KY������ �V��Ƥm.T�r��i7k���תV|��O���{R���\�@�8��R&���EA{ �.�,�F&�W�-��=��V����*�����+6qn<9?���~����c���Ʒ� �G�G�EA
��
(�ʊ���*'��M&;YFz��?�nˡ?�}�_�Ư)Rw���G�MA�-�(K�Bo���N��_��/^}MX-���/&�_����`�!8"�j�U��Gɒ��
.º�3a�\����� {�ڏ�������kP�/`;9G��sm�h?J-Z�Y(C�z*�ԣ�
]�=4x����A�����	�215ge���H-��\�9�[�jO-?�JzX>>捖���s�w̻e8����{��S�?D�C>=2�唯/�:����A_DS�M ��eF���2쬠eL��a�����]xc-���Xdm��lrQ�4�T�J�#H��.3�Qrd��o�\�ƥ���Z�"}��~�\�o��ԾY�bD��V�����]}�B��+v�ЃM�c���Ք����@����S��Z1�&A:�9�~T@�Yu��� �P6|��+�o�K��VRR�pUO׍���ݱ^#���s�_��Z
��Mr6�^6��~Ovv�͇�����O��֚4?1Bʽ���+5U�̏�����(`j�Z��9Z^2��D�<Ӟ!X��j��,/L����W��n?������"'s��oQ��T�E���Y���v��yR�a/ s�_��3-�?5���5$��+yV$+ą�|�.�
��5g�}R���O@ ��5@������%rv-�N�d��r��+':@[�̿�o$��I��ICs}L-�^L�;E+k�j�{L��z����f�as!����r�
,�RZ��uT�f��
[_�Il)P�I���y�B�H5Au4� s�>�@�K���"~wߓ�c���>�� OM�)�`�Ϯ-�Y9
�[!����aK&К�� �8� ��G�	9O��&4ƾL�JfD�W��J��5���ڈI.�~{v�MQG1��:�@�]/�Tuw&�#w9�)����l]��>�e�Bp�4e���[ox�r��r��톿�r��h����h�
���A�p�d�T�S9
���ߓ��U��� <�@��K�P�� �tq�p�!Mx�W`���K�x���+$JtSv��p�21�AwQ����7''�`���s-�4ȐӞ���N_	k����7�(|����*Nk��J/Ϸ��Q�W=:�]�����o�`�E����w���_���|�����sE�/�)x��KR_�⤎�M�([��@��΁����Pz�7�e|x��;�[����`�g8��^��j�#^e�v���7�$��R�K���\V2agC�<���G�4;D�����f�`��]V��:qXwgV5T�\�55��i��`t��F����`���������ﾎ��*9 �4V���N���^w��wrT����rK�~K���;]w��~]���I2�dϙU���Y��ȿ}����F3C3�����w�t�w{Nk��UV?G�妻e��d�X?��aς�*"�i�;jWo��
�I�P��I./M*�3PUefF)H�{�2�TT���]�'\1w���1���㇏_��RP~T������Jz��#�P����O7{�Qr{pm���7�X>�����wd�!�Sw��k:AbySS{�o���ћR^�H(����~����c�:�j-�E��,�p���r��ͯ�z�t���4��l�}��\Y�h<�� ZƉ�L��k�N!E)�l�K��I������?�z�7W�9>X����)�_-G6�hw�sf�j]�nɳ1�KT�З��~=P����ޛv�Y�3�,��,�&��Z��?��	%�i�}C��ۖw�	�̈<{ػJ�Z@��g��8�?_�[��1�avCL#z�,[B�U�G��4�^�|�h�鸋���C]��'��5�
hn�[������yt��Z�H�]>X�q�%V��p�9�T�(=�*��[��o���%�r9@k*Dt}5���f��[��7l���k:���Vd�^��aƐ��Ly���e���A�ٞ�e4����O�}��3��ϖ��M_B�gݠ�e��ry�r�c������l�o6�ׄ�UG��2F�� P��9�I�=[�'q[^�9N��}Ϩ����
e7ڛ�&F�,��Λ�	�<��;魪�ޢ պ[rq��+Z3籏�V���@=�&�mλ"��Y�D�<�����+�cfU	]�ː�Z��7[ �\o�d�׌gs!QG|碟z
�z��J���R�\���ZQ���@?�2�����23�9~Z�7��D�5Q+o�;���.��|#0��dϏ�)���k�58�}Lh�7�a��^�+�7X��	��}��*̘���%E{j��w����1�j���9V�~ӽ���A!V=IE2\+:���i��L躹��5�=��N1�:\����~$��x��K��Uf�]���+���~�k��"咱�34����Ɨk�����$��L ��U%�Tvf:q~!S�⺦s�B(X�:�nU�ܻ���%��]TܝbD|ۦ��&�E���&�墁�E3Ul�&���p"�78�: �^���VQ|�\`���O�Av���6*5t�O��1EBߥS^q�z�~���K}2|x�s!|�	��n�-��rwɏv�ʎޛ���<��\!�b���$FH|�@���s�Q�dαq��e�r�`��N�s>N�
�����l��^��ް* !���6nzM�>G�Y��{꘵�:��2�����^t�9y5���8����)�"�=د�O��@����S�����	/�:��^`�*�Nxb��ː�T�hَw���I���� ,X������ 3��.�l�ɟN�мe���[� !!����>:��4Ej2��j�px��� ���rq�rͤ�`I�����\{�-�n�E#�'�o����EύJ5`(�������)�[Ɯ7²|�������#��W�$�:���3z�D��ݡ%�!Ku�w)�w~�}]���9s�ʯ#D-�
��X?q`GC�7*+q>�B)�n�����$���$�sbLh�P �� s�Q�7�%�,�6�vV_|��6�w>O�o����a�3��.��!5֦��o'stp@��$�q�S:���!��p����t]�@��d�ޫ� ��H�7[���0CA��9�N�D��6����akL�jq�?���t68�tb&�7��W���m<}�'�����P�cB{F�Et_�c�>��u,p_���|�S=�[��sb\Z���c����7`Dsi����;\�s��i��:����Q,^�%D�eEWYi:6hhZ_Q�֘�G�:j����&E�Ġ��a�ŋ�/ro��s基V)�t	E��!�)O��M�\���p�:���	Fו���'
�x�@p�1x�*A�+�I��c$Y�#0�͟ݒ�����{�٭k �4����x�d�Yq�4���$q��pn�O�R.�oU�06["�.7�H�*��}�4��T?TCT�F]tx��5'\�:D^���)�0�H��/96�**�����3���s��Y�,9I�����G�!�̈́JWz�Q�H����>�
�TS��bp4@ Z�k!�����U-:�ne����,���1��$�؀�p��d"𦏴�L�[T���k��T�i����z@?����~��{�^��p;7�t��H;+�D�������l�[�(X�l��8���]ÂC��gA�@�3�Ȕ��\�s���=��G��7v�*`	vy�
��
)/��U�R�Du��͖j�Ư����z���	ae�hx��^"^]�f[���}�o��H�&����W�r���?c� ��qr<�h���zt����݅��*���L�g����^���y���7��b�ҵ�1� �p��/��A���W��]����Y��R�;��{*@e>Ȉ���}
b��F#����*�>.w��:��7�_�?ގ팡�Bl6�]�]�_�*x3.|qgX.^�Cx�򌁴��!"������}��}hP� �m�˯�Z:��r Q��~�ݭw=:j��#�o�g��[YFw�b?Z�R�g��{��j�!v��=�7�����&��}�{�1p�E8���6n*�i�y[��-������r©d���m�Kˏ;z�����A$	nA^���ū���M\#������pNQ��C:�}�~<� BC2�VUpfy�U���YwR�rH%uMٮ����48��z	��H�׈wB���,ť4q�9�T���A�}�s����l�_�'���q$����U�Y��"��Qf�v�ZT������nF�Wg�6�ƶ�<"�	�>HB�NMl��S'�ϗ�	fqX�Lޱ������x�c|�w#ls-'�mc��G隿��ʺ��%"g^SL�ߴ���6"=���]Ϲ���s�3�f5@����^x'�^!x���)��<T+���i~�j}�i^���';]� �w)K'�H���F��i�1��R����"+H�p��]yxK�%Vg����f^u+��N6�2�e�?d�tR �Z��4lVk��J�[ƝG|�>��Í�
�4tDmN����F@����ߍ��Ձ"���A����R���[ < �U{�L;K�«�:=�����+��xʼ��S^4m/ZiCٙ�F*Ȑ4��J�<�Sy��-�q����g�*j�?�����|�y��.�|�A�0�ZeS�33�QQ�F�=���<�����s+�g�/�ޗ��s�s��~_.)9E���Å��N��sz��5�H��j����	�;N���KY��C�(�)�:�:>xc�ص�0^����s�b��<%�_;0���"���-tr�|n�W��+�7~�$q50�mu�'9��x\<���
�\%|k�氅L˫�؁f�M�-G��o<x����l��k�}���Mk� �&�ή����-��G��Λ!�sp�d����O��]됁P��TMT��9=K�n�)�{Z�6D?SС7��+h˳�bdg�K*,�T�>3ثg�k�[�֔��o�c%b)�g���f���T��8�u��+NSe�0��e�=�����x�5cl���(��r�2~'�Q"h�A�sg��@Ǖq�hs���㲶���Z�L3�o-ֺ�=�ͮlr�ݗrf���C�ٗ�\a{z�"��h��G�������^%��݊�i�G�;'[����ζW���2]� ��r�L�A7z��=����deA��	��@���DX�E�5~)�&����R��u�+?-6MG�E���W�-���x�C�T
�TȦ��SҮSf��|��eTH�c���])��$Z�> J�Z~<��w�n~��.,��Lc&`	�#�˾j<$X�k78GI6jF����n��D�<*��!��wv}�$��)m�����m��Mc�&:�$7=�Et-�b�1=<�y�o�o���Uƺ&�V/����!�Yo��^���p�o�AYb���"��u�U��d�;B�J@F����B�㍬J�F����qȕ*����� ��:@��.拎hѓi	��� ��}�_/�l:����/���;����@N����*���߹��kEL��W��zdɍ����L"ާ��I��> �Q6,r���<�N�ކ���֘4�j6|��ljW�R�.�d#+�WJ�e�_��L9��nq���REG�y�x���AT�K������;޿*Y5s
*zL:45��d��R~���E��º>�SCY�<p�%���k>P^z��
.a�S�R��J��; ��xF��&_�@9E�����2�~�%�P�k�K�W-E��|�Q����Pd>HT��Pv�9��g��T���m4N�QQ.WL-�M.k0�g=��XCk2�>c)L0� ��_.�Dl�p�`OL��� ��-��Q���[�p������17%d?�fd⿪�:��U�ye�`ğ���P��i5UU�[JT�I/J���¥Cz�h=���ߕw��n�ƎM* i�؀`�"uL��-�-U�cl1�x��R@��-����c�@f%I�u����W���Ų����晞��p�^}��o�1���ͲT_}e�#�ܨq�Y���^9�b�3fŁ�,���q��X��)�@���B��Z֕�aѐ�F���O�k��(���XX>�Z��ڤV}Iʲ�𙆊��{U�{��k=��,�7�/ ��I�����g� ���A�VA"G����agd�λ�P~��4{����:j7�`,����|P��k(�;�T � ��� �Af5�cWF�Aw4�|;�n�e�֟��}�4�h����������ye)9Ջ>dl1�B����5�8����3��*?�����x�c�-ݼu�d������M�J��E�̷K�:��یRK�z�6J�Z><w�<<���o�W����[�fu�E��u�z��!����p���a�뒡eͩg�1r3y���Ke���W��$�/�rQ��q.�nt�>�H��e�p���H���d��n�0_Wֳ�!!���ff��7d��T��T�!ƿZ6��uv��ު"�[����l�c��r��[��r�n�j2r���Ϥ�@,K$��v4�{�0r�X^&Ř�7��	�|�s���˜��ʪAu,��m�&f�-���۶��� ���S�m��Y�܅.�#E�y��>�Z�^��M��(-��6G��Ƹ�')W�/Z:�, ��)��/\Ю _���u�D��OsƎr�T�q1�c�73߄�g�2/��<�����,޼mT������RafU|ck%Qt�B��������Y��5?C�W\Z�;�w
im�;��W���������6���W�>3L꡿H�-��{KɃ���$���5X�F`q<~�yË��c�����k��� VY9��h��sn^���7 طDv�7���FG���n�D�i8��o���TR�O��M��w��^��w~n��! s��Q	������F�I>\�?��ɦ^���%��k��	 w�8�־s���^��7c�����CJ�.��r��5�L��3���O[�>�26���Ƙ~�O �<S�I8�l�`'�y=X���Ҫ�{G��Z�~~�m
Q�t#��0��Vڢ�?�/�9�̈�oKi�,�p���b�$��N��	�T	���,�yw�i�kH�J��թ��s0���5�w���~��WK�(�'GZ��#�"〰�d��l�y_�Y6+C�'�̫E5��4�|�>Ce����fcC �������P���M*_�_$r"z����X��}�����i.y��N|���X;ȀL��7"�DwVM��Q^�AN*j��̭��ʓ��e�jqH�m�֝"I���Ow%��O��� �8���s�����Y"�������fUh��-<-!!:C��!:W8���Z�����6��W�?�;���2���H��/w�&�0�B���`*
Ť�-�:�����_�KFJ�/�8UC	siy�P�i�.��^�훖�/_�����0H�A�/"��	��lǱ$�B�4�nw�дn�c�m��-D�x��I�n�h*���{�x�<<7���:v��mk��^Mld�E�	��Ye��ɧ���X����}r[ꈗ8�RTˑ��E]R.Z�M1۟�4�S�C|�$C�µ$;tR�c6Q�	
��@�MFj�v��+��>��e�4�����o�&�k{�/f$�����R��~��	�K�[X���i�<jH�!q��N���7�:���W$�g-�1��<7'�x����*����R�Ɩ�v7��!���nV��`[/I�c:f%��VW�%a(m�Z�8�#l)���b�Eb(W��л�~AbjE�D�"/�1���.���N�\��}�#)�ϭ�����������V}.��?�+�ۡa餸���S֤��ڦ�b(k^�[����f���S��4����,�	=�o��yϋ�}�q=���ݷh5>U^켌Y��]����c:ж..��@c陋P}"GVk[e�i!&�6_�_1	M`g1���
�6��Y���M �Y��{�� �c���F��.I�F&V�	��)@��$�̎��d_�ϔ�%Kq��]l�n#�L��(j�m}:~P��������T���T�5��`s,�X[�<o��ݹ�Ͷ��90y3l�k7��/W�Q��0>�S��T��#�&���D.8BUo�����~�q�_Nl��r�K��Qtuv�i�4�1Xm@�� ��0�k�gP��O�8�4spM�� �r�։<����Cm%S-�a��{�|�	��OX�v���{բ���Wf�t�A�9q���r1���'���\r�EO�T��TCf����D�{YC��hRz�tLFw��n��S+�<5V)���4� X�6W��*����W��B�z�T*4��|h�BO�Ke����"3�w�
���m��?k�^�$8 �N1�U0�/�c+�,|��c�O��ý�����"ٯsQ�|e�ËD2�7m�*��*J��&s�Mwźљ�vTȲ�����޳J �߀����hH:���ټi�aP^�B�l�F���9��&톾㶂����	��9�Z��ml�뭶�|���0gk���Ƶ7(�E��h1��娯H��mq�g+F���)�Ⱥa>{��L�`*9�k\-���q[z�@��%t?��}�KRoN��\���#a�r�\��p0�F�`��H��绸����t/�>�%�^�I}�� �S��7�����q~�¶b�"��,���~�:2 �k����w��L�&�6�>r�(���,I&��Ȓ��M�A#���(~W*�V���R�WITE�0 ����$�5�J���6r�Ep�n��%�b���t��P���60��qa4�s+��U��A!���]��r�,�=
��8���Ơ�vo3a��6ez���� h�(�P�em��8�<���Uޟ�%ǆ��M?�u���w=�2C��f�|�>����%
gJ�{v��� ��v����C'�6�Z7+/����
�X9�D��u�w�^���l��f/��B6���)�Nkl9������Y:�ΙK.=|%b�RD��p1��ﶬt(a�S���\�iHK��ĖZ���{���i��DFy�]mC��(��Q�� �!c	K'ξ}v�/���]�X��aC�tE�����+���4� K� �F��0 ���p��O����))"2�N7l�0oϕE5��w�d+�R��16�aK鳘f
Y f4�AEA	��]2�	Чp��V�'�)�Jʡ��Q����^�(?�>+�2��_�;�a����\|���.�k�4���\M�dbr{<O�7��P���k�L���]�zc�e/�8��Z
&go�7H�`��B�t�B;ػg�@������i#5��J��^ ����b��B�U�ّ���u傱i�C~3���z��
9�;���?���
�v�_�6�>oQ.zK.��k5M��i(�߄����7z	��������	/�k�w��8<f��c�+ e�\�m��)+l<�̏*�g�40T��.* 1'B�m+ ���W���>3X
Ҷ_H't��Y5�G�����>ٟ�����+����ၾvr����Ĥ�9�A��O�v�v��po�Z䧍U^')�O|@���Its>ޝ��\N��� 1S�|+�i03�T��\������LI�f��KVf�K��K��]a0!�C�bd���!pb��p���lȁEȲ]�/ѡ��(f�)T��L��y��M��nQ[�.�� �o�B�C��Aw���0RQUU��	PO�W�gj�n� 92��#�~?M�O�$OY�|��
f��:s0��C�x�b��mnQ *A���p����P��Z_������TЋ��j�[:L|�⏒�F�QQ�Y7���>>�/���!�_���hhv������oWu��k_�L�jrZqڴk�9�\�2T�+�.�v��jG��h|M*���Md1��v��9�[�x)��B��u�td6��� �����|�s>���n�C�V6�����5,�O��q+�Lg;���K����³�n�۲W�9����hv^b�ųڍ��͡>���@�F��D�������[�[d��[��mh��憦�/S��ͩ�����23x�{�D��k3��H��\��|+�6���Ý۶x��~��wC�B��d��q?G��������Ӌ���\,����x½������Pu��l��o���T?����ٍHC;*����t��[��� �O��f��r6�(��Qf7�oN��v�s���U?H���[�[>++?-$�8f{����B1�B��0.١bJ��xF�s��}��tá����|�C�o�:/��������J2�6d��΂��ꆱ��֞;���Q^q�gdq�箋}��@�r(�oS��\<�`����Z��(�Y��-u������B� 1����0��S�o�M��,jU��:����#�jV�%��YL��ߕ�R��)��ۦ���֜�M[[�QJK�*�yֽ����?1 �4�ϧ��z2A_�pP��ɩ�i#q�`M��7o�+w�_��Ov֩w,(�o���}�v�mS^Yy�Ff�G
p����0G���Ƞl{�3=9�Л�y�r�i5XyB�j�y1-�w�ך�w�-��&�]J��o�-�wN�~�<E8�ᶍg�`4�?<Kk�c ��J���>t�9/�afo�.��أ-7D�l��H}#[�T$mb@�Jʔ�z������\L�k"�Qc~�m_�/ᙧ������$\'z���Mrx냄?��<! ���\LvߘC�v q�v`���ȩ�z⩲l�ޤ��'�>��q����u?u��p��@cæS@��ޭ{�@|}�",%%͞���8�;	o��7	ݡ5�R��6��p=,4��A����z��:���v��nۿ�X9\U6q֣�P����C��-������x��莴\rۃ<��?��>�G��~Ҙ����h5@��H05#dwuNد�6`�T5�_�}�ۧr]�h��\��S�K�6+�(��-��_0^q�Gm�".����g���7��z ?���(�G��eU���4�#�]{U������t���m�_���¯6DE*���,.�j>=P�NH���	�_�����K�����t
w����穼E��1ވ ���̷�:Ρq50�w4�;��qISb���E�j�#ߴ��ڣ�����׆��ARf֐\w�jm�+�����Cɿ��WWS�h�1nq)�<2�hop�ֻn��CzB��P.f�Y���5�:fx����|�%�Hǘ��Ø� �5�[<O��><�;j���M8A)B���p7���k����H�a��)��6�_�j7�~����EG���~�E�m��Uw�~��x���1b驨�b(�#��#M�_e7�����c�& ��[ڎ�4��]X퉩&���󿒹ZӐ��\B�a"�X��.���_#|��f,� ��H����D9�V=�ت�7IqӞ�x����F��}��Lj'�M�繯/��K	�
ܡ�?- �z(�i�e��V�1�D�+�꺉�A��vJ;o�X�9�Y�)�9��P����KB��+�Q7�vS>��#�z�\�n����^X��cl�32��>:l��<?��C�iG6g���\"� ����=S&p��/�BsM�50��΂����(o� �/-����Y9���DFG�����t�ܐ�j��ZU\Im�[�O?\9R�ȑ%�3���g�HR�9�F�裩�n2�����Q�و#�� c�j����YFؐܯ�s��I�4L�
�d ����|$~��=qd���ڵ�j�_:�0�1�����E����#��˛aƤ�#t�27L;�R�۸]s�u<��im
:@�	s8,Z�e�<R���_��'��p��2�����9��G���OVE�����?��J������v:���`ek�;4���r�H��w����u���~@�V�CAE=��ܞ����߻G�;)�=OO�?�$ ���Uj�]J�����UD��޳(�s�U���2��_B-qq�{��e�n{{b�1���YV��yy�&���G����?�
�ߎ�|#ؚ�U��(�G��h�R��9M$ BBtN��~!`�oN�����w}��Ů��(�w9��4T�:YaP��y� ���`j�RUV3b��ʲz�,JQ�??n��S����­���D���ovV�F�.�X��a��U�kr�G鄟ͨ:����v*�}����ڔ؇��T��H��ާ�������e��/�U5��z�I�����4T��V�����Y�}[�����
�8Hq��t3_j�eS�p(kTҹ/ۥ���V��E�,�6����<5�?W�C�V��R��xBݳ���?�1���r/5��5m$G�$�C}�z p@����	ģQ͂�Y��e뚂$W�1����9V�4d&�[���1��*(��|�q2��	�?�.��ro��y5d��[^�_)���`��L�τ�Z�%�Qe���5,��Z�>��W#��]��ZJ�ĻF��=d��� 4Q��v��Q�ƍy�����d�h-�y�/.�����lD�d���;��1�l_>|Cg~9��_�$z�F����i"<5ݢx�N �G�8�e�<�d�S��d#�"��[�lnGJ��V���`������2{M�{�[v��-��/���h�8S�#_��P�*���rt>li=��m$���� ���{�c�Ly�H=���y��,D�������`�T&n��ݤ��� ��H�-UU�g���0���ܵ�>����Ӄ��_W��i:����k ����.�T���ƭ7����6j��|X��Y$���<��v�o�'z�Tl��\�vF�Wp�E(�p��/���dX�b��;���[K��^۽���x>ifW��BG����ӚM6��h25��(Ա�{\?�;��\�o���;��4f]�!Ke
Շj�=�˅?��ZK���?�+��)�9�7����ßM�'N���ܵ~���;�t3�0�JTl�n#�n�~W�� j����b���⒜3���Ӄ���@js��&\�D:i҈���DL���K�Ѐ�6��-����e2�w��(�����]A����[0K��7�~ǽ���@�j�(m������M�z,�Sq�#��K�Q���N�ɐx���UVS?
j�k�Ԩea�w�{4A>���5v��Q��TeĀn'��Z����N~�۶�˙
 �S9��M̝����P�KT���Sc�߱Ё��EV|���c(����ؿU\�����6Ã$�u`=	S4�}��j?oA���|��[ܰy�JIq\�ҖI���S���8i���$��`���Qj���ci@��2��y]=ܸ�߅ߗ�M-+����`�0Ǹ�3P7�j|ox�{V��i���Z1�	�Mg�X�<�}�� \!������c9	���s36��K��j� مw��$�5C��/�wq]�kpF��vK4��m��a(�8�G���.LRFuH~~��&��r�<���2���1�Ԕ<̟0��|����\��)�ln�Z�%y���|gۚΞwu�DPibڕG��A��r�7C���S���q���CKgo�.��^	VS�7�O��;�G�q&�c#��9��/1ls�8���
4��Y�?	ԟ[l�P��_�dY2d$AR�6�H�V����lZ
-L��ts35����#?����O
����"��D�t�<��+x�X�16�uչi�k�Vl��j*2�E�Ri�M�O�h�F�qr�A�djу򏉽����b�����)D��9#����d������v�Jzm[S|_O���Bfw�$t j6@�� � CLu
C�H�	�P�K��'���x���"��r(H���?�ȴ�CeNe��&�g���p�m��%V�2^SLR�F�C�����g���>�73��x��9/Ԋ�=I����΍������g��*�������?�#5�����v�Q>����̸�7o����&<al�v�m閿?�qMt7|Y�8��8Q��w��ݓ��ƃX\V���cө�ЉE�X�}^,VS�d����)�Ǳ��eŝ9��6Α��p@�V�m<��Xsw�Y������?e	�7U�,Bt]vJ�X'�Z����t�ҝIJ���0��C��{�>
J�.~���O�|�3�8-��c�9��.����S���'`aOS/
���s���姒ʗH���>�>̞J�p���9�(�`,����5TP���8
�;`���Wo$�*N����Z�ř�ru����4u��̡�[cu�!��O�en�s�_O��k��#>������5��]���3Y���A��N�ݥ�>��nz���p�<��˳��y���a	���k���5�	Ѳ2�j��,�)�-yh����П��N�=>N0k�ߓO�)K������	]"9��IA�}���Paݚ��>B����e""9ի��ibA��L <�!r6�`��Xt�p9�C���0�}��C��`xq�w���BwI�G�@�u���؉D�-��5(���al�U;O���EoFn�f0�*\��(W{��vT�m��:�@3�B�sGyh����EղF�^N���|�~�6�;���(��[�Լy�{O:��*(��6j��\,�D��
"��}
bϲ����0�4���[���´��~Ic�����݌�	F�1iyd�ڸ�-�����Z�a���\��(����g�bϯ����Dn����CU��t�9e`h`VYŶ�x2<���`�O~KɿU*+i�F��(U�^ ��hQ��!W�����Ufިg��p���sUfi�b0����Q���Иy�%d�y��.`�>]�n�-FalS| ��Z�M�%
o�(cH�z��[b�\���\V��۶��{�C�6a�������'�Y,�a��Ӑ1��}-�$G�&�����V ������/T��4b 1h2�G�Ш�VnΊ3��8F�Z��,����b3e.��r{W_et�m�Z��)�O���5��P���*�غ�u�"P#mC\�E��T��[I'/��Z��`�$��4̘�_�
��W�K���o��Ǎ�c���2`{�������j�s��a�z�LL�r�eI�[�'�Q�p�gâ��B]��A�s�!�c˅�l�j�&≳.��6
��,�R��c��"���F�j@��b��4�;��}���OC���o;-�)d0��C�i�\$|+")������L�O���h`X��ej������ኚs�}%KES��(V��j3>F.-^ˀꯎl`��Wq���򯢉'�����٧Z[��ЅI�>�'�^#�x��xGiD��U���}LVf����M@�Z��^:���yO�=��}�W���Z�-�x��4�� 2�7E8seHײ<d Yˌ��d��i ρ�LxO�n@<��8?���:
پ}��4��+r�#X>�2<t����7�����R1� z w5֜�6`��js`�$�������]��w��z���]�U�REj9�p��o���mTu?7Sefj�K�<�1����v�q�U?�c���{�M�3�����҃ꢒ#�zA��W:�$ �3=�'��L��Cꢲ�l:�J��=�����l ܢ��Bl���KiT�bcvt8���ť^{W���͖�^��s��/o���*6uR��F�ێK� �Ɉ�&��5� ��sȿ��C�y���/<�3d�ym�m���I{%A��C�o�Z��/&?˹"%�M9
&���=�o2�9��]Q�D��H�p0��K@�-,�v���t �1V�x~{�b�?/�����Ռ5*7�� ��yx��ob)0�?I,ϙ	�}PN^�������Y�? N��+�=���~axih.��ޛ�N�������ߗ�ཀྵ`�c�F'�O���.@�S+C�L�^2��y��^4y.�濗�|ng��3�s
D��ݛ"+�[�I\)m0T~28~�ơ�%8�0e5�L�t�i���k�>�2�v]<*9�O���B��[ޮ��YYM6��c��X�ӈ���ehVzV%(I�j�S����"
�m�u���EG<[)��Y��/D.9��+	Zվ�z��8��VA���I�pbx�c���&��'��I��pF�~���ؠA-�O���~7�ʔ%G����w�r�f*�@DkAj���o!,� W���E�]\w�'}br�KOR�wx���,y�HͲg��^�H)om���d�9�V�w*v��u=%��%��?jG��Q'J0\nK[w�����,Y�ev��K�t�]�Ue��M��b�0�:b-$*�V��
^ߌ��=�~�s�Ji��`�B���s_��G��t<E�ƪ8��hTgH斎3b�K���)��Dx���ϿE�[�k������S���� ������"�$������Ѱ*�}��c�ޣ�d��g6��ގQ�̃c#۱�:���Q���|����꺺�x�{<����>�RzY���)$^����ڲ���=����?.Ѩ<@>��&KS����,�r�E������ZϽ��8������I�����מxx_��I����묇wt3#�)�^|��SS��UfP/���b�a���)����[��]c��f�$��QU&Y���g�Z�2��?W�����C0�|b����-�F�b��v�.���;B�}��B`����M��qԵ�GB�\z#�A���Z���n��������d���{ށ�ɉ�gEY�X�3~�U'��]�B̷��02���^�!J�e�!���$�؍�t���3�4���oZ�ܶ�p�"�����h  ~��g�L�N������Q�_��&��ҩ?mB ,&Uw�z%���N��z������=��G��Ї���!��/�d�3Z�����(��⻆�pnTjgx�M�g�Ԍ�G 9Kf寯����d�w��]�ď����%��	�~}(R���8CzZfꃇ&�[�y�А��{s�5������R����A�0>�@ඪW|��W�C5�ӊ�u��qg�?R�*�r������K�U�M��ݴ��ۆt�������lq�������>��e"�>x�s(�p�9L�Q5aP�s��Zp:j%55v�@MA�oS#S	+,�������!g��%{�8�Ѥ��a6���g;6}�f�ǜ����w����$Q�%z� �|,F&-��N��[_���x�V��>)\D0\=���qc�X���]k¬���koܦc͋������A�$�A��/�ʍ�A�p�.T����?HZ5��3}�`{�\��S��cD�س��V�Ȑ�Od�i��tm�6�ک�w�����x�ӝ96�7�]ϰ/���LHi����0'i�VF�O�R`l����ī�8�ٸ�[����6����� ��
�f�$,Ѯ�����)ٙ�J��s]->3���N��x�k��
�x�IJZvj�T�N˄ks�PL3��Kr�3}�	�L ��F��ܶg����sÀ�lS�g�	!{R� R�(�Аʛ�m�B;�-�"�\�<����;B��<�̙�y
O��Z%�sq�C��@j��v�h�G���sh`ǧ�Qo�} ��hC��3���.���a�E/��S���m%_��ҒW�E�J��|�r�W���~�-�5{��PnX*��e]4P�����>"���Ɇ�1�١�ⲝ�ӕfa<���O�w��"�%|���;��T���!��P�O�~	Q��m�,����,�%&�+Ŝ�=��5�[/��S�$^Zqr�B�1-�s�)��o���z��HR�<��K
�p�3¥��n`�ȫoY���>��,�K�Æ��f�D���l�c���x�����ip�� ;�����"�M9�#�����k�/��d%>�^N�J����\ hψ��X��)�vVP�*�3Vpk���E�U�e���L�x��d�ȃZm�#mn��[źg�G0�j{��41���� 㬫��ҧ0 �De�J��@�&�r(�I���,�D�v+A���~岉,�⾂]���(?Y_P�ޥ��DU[�Ǿ�?�8���t�>�6LLJ5N��^��s�"6O��1(h��#OJ%����\���-����� B�@����έ_��0=��u�i$�t��o��v7�o���L�Ya��i�uR���Y��ӎr8�twW�a*���-ҭ����V��5>����u�}�V#�h�k�#ؔ�ݬ;��T�ֿ�����3Yz(���;���`\w.ܾcg��ߟE쫖�\F&Ju�Y�x�Xm�+,b�5dGs�����Im.Bt�n�n^(P��?�%Dr�e�#J�ST4}Z��H�Y?G{�b�4�>ǝa�'��m���B`����G�m�սbc�T���|�4�*v(+6G�͉;��1z�v&$B%O��/���[r:��w�d(�"� �s�(���a@�ϝ^�~I�ĩ������貈�bl.y}�s�y�v�𖏫�ק�Av�G���2,��X]��S��+;~�f#q��J)0=c��xt����խ��JQ�灜f����"S�_�nHvGd���<��/�L1蘫0  Ț��&�����ö�7��U7@�!Ar��y��n��Q2���U� �/���
j�b��k|?�0i4��0ea鏥���I��v�~0�� P�U���'�EP�N���??\f���U�m�>������'_J�%� �g��dHQ�Bdf�h�)YY�k�x&L����
�Y�~�L�TBs�h_�>T���k�o�hvH`h9�W�z���̡��i��Z�6�e��Yɛ���0Y�CA���e䥡�f�a1UuK1�EnB|H�$<��ɪIc�g�}(>W�<@o�E�m�z}�|��Uu��-r��{y�L��ܿ�)�7\����%iU��Z��@��4���A���/�Yu�JW�9�W�ˑW��,4������]��u���N��lcZ�L��J���%1\^�mb�q�
�qY"�DT|&�i��GC���2�C��}�^�rZ�e�6;�x�?Y����Č^�-t4 ������ۂ��e�w>s���Ą��2쑽R����`���O��J��7�Q�	he�~�4)/&�s���ܓt/�����Ç�;�l�}:�9YG������m����Pݷ�t�W��͟�l
`_��Л)9P�O�x7�' 6�����u�tJ��35�<�*��V��x[������O<n��3*�:!��>�@ą�X��>R�<��� I�~~�3a'B٤����f�*�-����&7ٝl{
��=��1O��*̴��@Z�c.v*^җ��\�����x0|i�=aX�V�*�W�{�H��Q��K=X��W�ҧ���������� �ci���ت�瘙��6����H( 
7��OW����Z[��?��>�ҷ�l��Z^��v%X���Cji:��0Q��Ă	RK�Y�{� �"T� Z�Q05k>Wp[^b��.N��^�;��,�O�T�]��0M�x_�8��z���i��P��f��޸� H0:Z@ʹ��/��!�1]��@�Gd�G�Y1��j�k�tЦȦh�C��@���W%��Q8�:���<����~u�n�铰��"|�����VnB &�T��@S�F�Qɕ���v�ꫭ�y�*�����Q/�4H_�~0�<J��r3�)�{�}=�~�����Ͳ�c�?�qZ�U?æ4Q�ڏ�蔋x���2i/�?�y�[���1϶N��9M����;���D���~�-�˸�`���CJXJ�S��ǹ�o�iz�i �p+��>��T��<���Ia�}��;J�N�_	8�������Ɋ���������l$�,X�̞�����ˍ*�MM�Q��3� �I��'��ܭZ�qם8�XlFy0G�0�ְ�z�H� �SF��Ѫ��я;����\��5=�ϝh�� ,˴��L�0�����,x1t� `���6�M
����X9ؤ�
Z���vim�Da`M�%��.pt��f�D������vx��~>5e�TF�g���6N�����fu���<s���@ZL�X��G`�f��8��MA�J�y7�̤�Y
G{+
�wS�[:���O��f������������@$l�h��N�I+��UJ�c�9�p� ����`��^�%o���"���_����̮#Op����<\Yt�@s�w�U�Z��Jy����J)U޹��uŲ��P���l;���%��d�
�X�����_q�L�2�����@p�̃�R(i�dB�Y����@�D�ґ��0M�DS�-�=��'��!���T?]�5J7� 4�ìx�k�'��RR$��I����@��O?�&+��
A�
�Uux(�h�б�/v	t�g_˩^�)�Y��s+5�.Z ������T�(DG�M��׭�R�G�U�K<���Cp���%�u��pҤa[i2���w!+zMJ��%q����a�Щ7��GH�F���	E_P����|���F��j�!�����
ѳ}���5��# X�D�d�-���=��2bϓ5麺�9/�%��ӱ2'�y��M��}}�W��˷L����΍~�jg��,L��#<Q�4s�������r ���X��O�$�b�?��~�MdoC�S]?0u(�G����2���C�$U2�u�O�o��I��Ӂ�""N9����C�f_���
��OQ��&싫�)Ӆ��D���4��ʩk&6JQDVn��l�bCp�'X�^��(�o���/ӧ�w��'���,>���	=@�@��q�$n��q�� �_�8�P/�ՠu_��-��7�5�bC��9����R��|���s�F�?8l筵sLx��HP�w�$g�Z�G�E�B�/���r�Y��`��5d�b����7��$�x�)mq�8)�(Hk�x.-7��;�L~�֎���}@��CO�F���x<�����8S��l%NX=�O���H��U��n��a
�+�$ָ�j���r���u�.W?�-�w9CZ�雌\ô��K��
1G�h��Sƾ�k��:����,ˋ��Ȝ�W�gȉ T*���� ���J}|�V	4玧�S%�3�牒�X>ʢ��xW�������P�eV�eA��M�3�'aJ�5tk��F?�ȿ��Xe�l�X�\��������!V���:�,��Y{TN�pNm��{.�)�1�NQ꺓]n"v�����O�C�_��(��e�C7s�ؿ�@�Ye6v�c��$�JZ�~}Zp�g#��:#o&����n�B
L������:>��pX>����@;gv�'e)�h�ּy�e9o�6�L*J�Ɂ�B7A�	v|M��� �m��|���a@��S��rn#b�]�+;�:�9�Ĩ��:��=|݉X1
�
��=����Q4���S$���04��JP٢��7�B���_��Ru%0|��Y^[�fW�6�Ԉu��2;��qsw[m�E}�C]X?
O�nH�7��D�&���������8����~�0���f+�nEhݝ�~ēѧ��-�
��ھAOw���vq���2��׸���/?�� t��LI����Ce}ɜ��n��L[�x�����s���<|��<+��@�n�i���1*'�����������Z9(cU*䁲�t�?�J}��y����Vp-.K���_V�2p)`����8��f=|hr���?ŽފD(|�Y4���$�kZ��y���<���+��5e�CGY(Д�\�� \BՁfD�=t�N�r�v!-���/CC�i�Y�:(l�{z
�#�͍Ԍ��&E���Xn��/r�3�_��m�k�7���F	�S�竽IJ%�����t*�r�L�j���3n(����K�`I�R�:�����M<�����D��G�OI����N��z�U87����Zt%�B�j���4��� ��U�MI݋��5klq;	�8�<zð�6)�xT�ذŚ�����]��(��D�8�ީ{tp�ohT�������߭\�"�6�x�����YdB V�  n �`�[<�wj(�V˰C-���^�*v�Yｽ���$��ے�#-�Z�Z ���%�d���1�Y>ny}��L�B2^8N#�ݲ����#�LF�Ţ���k���jm;׼�nWj�G�N�GȎ5YTav=,D���<AI-�h �lPOR+��$�t�=P��oZN��xdO}g����71Lt��LHK�FR	�}p�ʼ@�x��=;��(U"�5����������Q��.pY��G�yh���"��0v�܂ ������qW��w0��~�*�s�L�/URQM�e�j��,U��3{�i������~5U�8N�� ��Ώ��wު���w/SG��L��̸��A`�@���=8B>��>�,4����+�HHY���3�����h�DK�Ь`4����/I�fwg"�%���c7$G�-�*r�%�J��;n��S�dBe) {,7����~r��DO-cæ���ΡEV���H/OK	���&x�΋Iz��#��WF�j'����#�ԏ=����#DI����40�O���F~L�����ao��=��H�˂<�@I��� -�"���T�mU��3'�:�=�ٍ]Y�Aע�b�g/�794Up��k11��X�����Ȗ�δ�G���`��u������S��jn������h@��@F�S�Á	6΢ܘ�j�m�4�ャ��N��9�@�5�l,�9���~
��9�D�f4�H��5ЫZ.3Y:L���4��h�� L��I��X��t���z#Cj@����%��mO�I2�V/�'x�.?���U$��W7�r�����9֤�Oñ2�^�Z��zlt�N��!m� �VA?���pyq����$*WEd��h�4�y�� ��<��4[�ǯ���E��:4���2�#����B��e���"e��p����( ��a����]N\l�ae���.p/�V�슽���E��!$������ʹ�;�-_�`	�?ڳ�����_*|}z<�b�~RB��<���k+��k�A���)b6�e30i�o�mV6�C�(��B)�*�W�rk*��`B)h���ɁX˫ c\i����MZ��JmU�DsA�:�7�V�A2��I�����_��t��}�y$V�:)�e�Ã3�l�3�Ӆ�r&K��.�)}_͊�����B+g��/{*�y�=���['�L\��Y��5��Țm�w�v֖��Щ���<B)E>���g��Q�M��LZ|z�M�,��Վ���w�m��5���sp`s�3mKP`��t/��`bq�l;yI����v��� i���^����(B�٩�Z6�	��wϵL V��v����׃��T� 9S*S�9�Iv�����N��~4 1qfT�e���_�6�<g�B�ѦVYB9�}�ަ ����9�!�e>{'�~޵j�2$
��w�o��M��!��I���q3�ȍ҂�����:�j���j��Z���U���*���G��z�$4���=Z~��Y��`5e�ٹ"AO��M%�=��6��v��5��WcC�m#������'�Ea:��@�QA`f4����֖bU	q���I�L��e�z'2D�m2�}wXCnmoj�L`���	�y%N��O�W&�T� ��<W$�znϡ���=�.�6�/.�~����Kf�+�c0t�S�"J�E��� 걝7�Ib2+#��-t(@���0=�< u�BV�_���Ҁ8� ����}�"�}�PoS���&J۵�[����f�D3���P�r ��1Wл�z�W��@��ؒ�=�q����u��m���(�(lQ�X%�R�&�Ŷ# l`f�U'���o���F���C���t�-�+馦��~2�?�Q���y�+,H���&��\���'�׹*����A�`�w(�<��;jQg��<-�X�Zl�����B��w����VPyөǎ&tT���}6�M�V�z$1��]��a$�Rr �崳��{*`����V�]**���?�W�q?}�KF|�%�~�����wn�"2k$v��87�Ĝ~}8R�&�4�ӱ���p�����yRe�>z&`/�������u�*�C�[&5�OB��@JH�K4�ܩ���o�\{��ؼ����וX�3�!Q����.p|�p�t�ْ1�xt��`��J4�B&A��
2^G<�����.���G�����&�4>kc�(�<?���S�vd�F'��#������2,��Fo�
]�H�x�PEePG<�g����&���������?L��A��.(H�5͊Y�S�g��P��9=���;y(Q�#�5�i��}5z	�Qe��AI�k�c9tyð8�xy��V�Sѻwp��[>r@��+��;����Ϛ�j�o�@M���_�����>o���'��rP����nt=���m�M;�A�I���_T{O�o��:��+�<��i� �iV���S�|�|��;��<��� �,tY�{σ�(�g��m����%���ŘFړ#��7�/?�pl8h��³��p��ޖl�� hҕ4�j^�<�77:�[��������c����$V@C�l���hX))i
�L(�}��*����}ي�nb��1�P-��ӳ�ڂ��x@���/�"\�]�SE���EZQh1	���� �@s+�3T��a��خ��g1\����pJ�G�!�b(���?4d��I��foKm�̬��I<]������~�E��K7W��k�F�
�Ҋ��;�b�ѓTy.m������;�K�����<��ƶQ�f���	IF6'����T���M������a�w37Y1����h���z#ջH�̛������F�h�\<��0� 1�.A�*�7���v�O��/���H=�B�M���JR���]{x�2�QTj����2^Q*���5H'�ơ48k��>�b�YO��Z`^�]([�h'�,����ʯh�)���<�����gc�0���7�bG�����{e(9y{dJ�z7�c�;7������;���s��M�ͮ�5��� ��4����V����i!Xj�m��fB��W��
_>��7YA�হ'i���-�q����,��P��V�a�V�E����><�V4F�Dރ*s�u�G��F`G5�/ 1�T�a�B���Y*g3��R=��!�~�U�_�N�9�̫]����e_<�bR����h����'DƔ��%g~W� �� �t��Q�9\j���wL�T�Ǣ����2���R�FZW'��*R��R����=*�Eqě]"��!�H�ɦ[mdm�Ǯl���\��<p�L��e�p ۄ4�jp<a�>��.I�r ^l/��\�2�>P61h��jh젇Gn�S}j����ф�5Y�#:���97l���<��% r�+�T� i�%��p&+���<��6�c�8E(L��y�| E*{<�ؗ:�@�Ȉ_;���9d֔t�mWũl��&a}���L�3���1M�m��ie������k�
��T谁�6j�H$_k���)l
�N�r�M�SبA�t�����豂�#�8���Cb����0R���D�#2����Q|ETAHي��� i�Kp�ߺbU�tZ}�D[*.� ����2kc���0~����6e\���h9��m;|F�`��;U���k���~�q�C¡�C��õ�� �m�;_��Ҭ���y�]2������=o]�����2.��dd�;��j�����B���d$y=�����wL�s�H��S`&~Fe=�е�M����ߑD|���?�X_2o4dԒ8ĭ��ˣ}�ۛ��`�TT\0�7������N�_=���~!����C�Z�F�7Y�+�����ݰ(��	������תIU�pCmJP�N��S���u��?ס^�۽�J>�������8S�Ċ��29xr�6���OZ���f
��'h�Dܾ��Ģ@��={G�`�h5+�l�ُ�)��2Xol���~6�"o�}q
��� ����*���x�>���' ���^��a쏾�zQ-����y�F�����ݯlt{�/.��J��.d�mGlq�_}��Ad98��.������Asz��-��t9����^o&&�(�Ѻ��K�MFgT��ߥ�XN֝�	�늍a6R�剫��J{)���9õ�q�T.�?�=CԶ��xωK��|���stk��.O�Ԡg����#�O�zWw���3O�:�5}�1����)���&�_=�3H;|� < r�]�Z}������,p�=����^�X���X�-�,�Lٳ�0���k��M�\��=��iz\s���O��c�N���*fs���������Y�[�7���Ɖ�؝��c���ۅ&o#��C������,V���w�2qU��DiO�fBv�LH{�R������U��v�����Z&bG��"m�����E $��S�X|{�� �4��m���(��
Y����UM�&XY�fӡ��ag�2Z:o�g��\@�2�c �2������CҬ[=�|�-��j���ғ��J,��/Q��C�4N��R�'x��jB0��P
�ނ����x��3R�<����O7A=pO��"�����_|ܞ�u���~L�����o߬�l������U�K<��Rs@lnT.F���ɠNq"jE��W>�Q�Z�1u+J� �Xb��y�x�s��AM`�s}^��̶�覭MP��k�8��f��}��$H����������f+��tt�N��G������:F|�I����m���\�t]&D�f��+�FymD[�v=�nQ���خ���b�-�S���W?w�{��@z�O�B�fs��D��^����r-�������,7����L�?�DM|K�
�Z�_s��g��/���_۝xo���u}w&S���ŋc:���e��箤�9�ĈR�s#~��*;��#^E�*�K�Y���L�l��JFo�.��t�H�X��'N��Ĥ�ũ��GV�6�n���;N'��v갹=+��R����]N���t��źeR�������~�O#�7��|-+���ͱ$�������t\���&(�|�XG~��-25=�ć�	����5{�8��<iW�B�4���u4��N@ٞ�,Ь�P��!#����^y��-�Th�Z~���؊:�X�t���0ηKNB����	��c���e��_-$Ұ�JA�P���ftY����s`��9���X����K�Q(�In.>�Q_*����	4POڜ�Gm���yܵsܵ'���ͱ9��sm�l.�C3�"K�ܳ�|�a�p�l�q�NV�l#�x�'�k�N�U����W��~7�����������궊�Y#����V��͞ݒ��FȚ��L^&�:�I�u��f�����r�t\�k��K7����D���2�j+݇ޗ�<KJE��9Ni��G	��V�FD�Y��:>��ɝ��MT�EA��ʋ(j�W�XU;���q�)�Gn�&(K�ţ�]�2J�b�
�"Pݬ~�l�w�Z�Ҥ_�6"��emyN
c��������{p�Uf\a�-�^L�L���s���&_�dƏ���*Mf�j\��7�8�k[������%�'��d��KS�n^�G��4��46��J����a�7f��(pp�ݥ�H�N�.�e��lue!\k����D���Hd���{��z��X�h�8�R�i�5��N��iև�m���W�UL�[-5t�b���GwX`W��楇}��V��Ok���r�0`c%�j���|5�_��@�X_��c��A�4��n��}G���ކZ�s���nw�ۓ��f羙��j}��j���1�J�ʳ��]�	���*���PF����k۾��ηC�Z�x��}�Iv-�S'�(������߷`���V��P�$m���L�S�v�ǧ�̡D0݇��n~���xR��˲�������ֵt���u��^֛�a�\��N_�)<�m��ʠkMK��0��>l9���$@������,���s�N!�����+${(���M�JJ���ύ$π��3����6�8���s����P�O�%������������ґ�����GIИ����P��k}�A�\�M�e1�n����{!��<�q�&�	7�3.�MT�:�:0KI�]��YARv�ضZBHm�.�.!� M�l��������)�Dx��<�0���VS=a�����<P��}.V�ؽ��������i��ڗ���w���_�� ���$O-ϐO���0`Fv�����dl��֞��1Ǻ&rE�E'5��/߃�$��O��[�
��Y�3l����	}�VL]���DF�O����Ӈ[��0h�L�OI"�p���'�M�ׂ�C=��C�(�X�n/�)��v3J�d���C$\�E�;���;�ݧNd��^.x�N=t}�3�NziJJ�̎��mk��"�eπ��)/��Fh�E�4V�� |����g���z�-\4���I���:�)�(,�ìSS�ؾ{ @�d-���y�T�|������#�u1�	������R��x���nQ=3�㺞ݗ���J��I�����lȖzT�[���j_(��/�W;��E�ʞ�-�گ`T��T�o7��1�c���REGU*��U�6��%H|d8��K8+U���B��w�?�̹�v;1
b�$�30�W�|+�~8��Rs��暣��Ӗ#s�'��:��z=�阐7�Bк����x���aBI�/���a�kv��e�x� ���*=[�X2��ի����J���O'�I�E�b6��*hA9����n�!��5�t�Y:�Hke�NЮ9��n|Ju��"�F���(��1�������0�۽}��&W�ɿ������{��o}����ٛ5I��\6�I�(1��S';��u��"�ź�3Y�-�5�� �+?X:�b��(b����^���}B�2�2�0H�'^/[%2=��b-_�G�0mQ��A��9O�>���D.]]nԼH��U���H�
=��n���V������t<����#¥��E�>_h������I�娍�_4��WI@Z���#��D��?���&?�~x{��Np/�A�x�.���w���ʜ�9��/$��VSP�� ���s(��hg<Y=�ZFԿ�S�|卟R믪�8=+��C^�M��������Q�,��г}����;���>`�����ln_�ji֍��h�@	
Z���LT���ڎ|���Ҳ�DF�_�TY����Y?e1[���#_���S.�<��L�FS�UG�Z��d"W�t�ָ���Z�=���V�e��������~�z��aj���:�G�y�����32,�Cp��Ǵ&�z���XUo Si�»aC�y����.�z,����k�e���5�,��bh�:�i�SK�/ޭ(����uuD_s���Г�?���"+x���-[���5�Ѻ��y�C��Q���[�|q��Cl� I�\�2�����������z�?
���)q�N��܍3�Q����=_7�UrS�|��u��$�%!�h�Ry�k!C��u�K�����x�g����u6>kMݐ��ɹk��Y�b�mo�k�%��/ �/_��/K���{!Z/,��9f���Y=�u���l@��	�����M¡����sbA�s;���O��?K�J��HK+�u8��b�N��$��qޡ��;�ʇ
[i\�;V�N���>�Q>7�T�A��@$��&�\q~ѡ�>`�Y������^�A���d���:�����|�?.�҆u��l�d���=1�V�dB����w=��y��D�s�5:H��_`(c�?6��C;h�D�6mQ%?�3��8��)M��91��q5l[��)���b�5P��;�-�a��[iLdm�z�@H35��@vy�~�^��?���@أa?��d�=�a:Bpdڱ�ii���Ndpua�M;AcJbC�p�Rx� ���~@-?�Ψ���X��o'9g���,���Q9�_��[s����vئ&�b�'p��Ga����W����fx�y3�jP�&Q���F�f��f�Y�2A!�a��|�|ˋ.3���Lz�V��qfT&&�h������{�r�#l��;(������и@�
��x}:�)�tk���p ٗ5�|��z�+���_,��\�ܟ�����9�PUe��j[䱼�Q�T6��孨���LH���a���!�������E����v�6*�fn��gC�ã�%Α���P{�ר�<ڝe�+=��K?в�:�E�Ƚ�{���ds�G��)�E���K��g ����H�X�
E�T�b�S��!����K��RRU����4'�T��d>���mJtg,�Õ�ذ�*��_i]nʉ���N
7��M����0'�u��͓���N,�d��n� K9 ��W�� ����RoX:R͙o�*�?h
��}y�-�b/�Qr2<��=�[��KR�֩7�g[q��qY���GK��D��(�O���.؆ U�2>93��������j��t��]�!o����g����:0(5��U���}��;�{�Iz6�g�J �+�-K���� ��WB�B̏#ߝn%�UI~�:�pR�r"�1La����HZ�s�a�ǳ
h�zv�o)��6Ð��pA��z��\���:��H��+�V^i�a��U��iu5h\M#V��>��#v�\���h��E�����Z qF n����������v��S[���3��ೌ���5��ڮ�w�4�4[
�Ë��.s_�m���iz��t��yg�g�q���ˁ�	���IC;KϮp��}p������W=g=		�t2������k!��#��8Oe�ݼE	R'�A�Y&�{ 6.�-c���?��1|��!�{�����ؽI����OO�1��UK���4��B���V�q����P�zo������*�'�j��/d����tS�� ��?����R��V�{�)���<�|�\Ͽ%/���s��k���+�������S��?5LR��MH,Vڼ����V������k��J��I~~�;���1.n����c?����O�V�_��zi��0w����e����J���v\���Ȉ�#�$�g�L���m��o�5Kr&|�����7$_%Z�)CVu���3�x;�>��K��a7��}YƝ���8��d>�x�y�6ުH�����8��0U���5�����1/�0�P����_��2� L�Y�E�	4���o�pKr�X�/x���B�dJ^Ux��x!򫀈R��G9�����hפ{V�H��r���S��u�z�a~����Ayy�q�9��"ߌ�^����������[�b��(`��AdUH_���i_CyJ�DeE;XW��ѧs���� ��[�8/s�ȷļ�����*�YA`����,t_s_��D��D��&>t�7jfx��I�� ��0@�@��v9���%��a^��/�,O)�K[����z1r�Ϩ�Q�j2C���+-Kw=SR��Rr|�ݵ�#^�����d�F��<�evE���"�{6׀!y`|:���w���y��I�h�c��M�D�@
��䄪Uk{ ��Ϩ�k���V��,�9	�_�a�y�/W6/m�4kW>��M,E�U���$d�,<��A��02Z`����\é'F�����
5�|��#	����:.��
Zh=*���l����P��)k�)�ҽ�f��ѕr�ʱIg�Rh�P����=�`LA�?�"-�{LDP.���]Ø�Ed/q"�����K�em��S�"���8	�ɽbP3����K
��aqO���4��?:����{Wڎ3��0�|IS������b��J� ��=���Ԝo���݄��g �/�0󃋰�!g%�4��Eh��;3�$��Ȥc�'��7u��#�ES�1T+~F��r�fh�O+��%���`�s��x�ŋ����� ����Nq�U��C�Bư�;��q�)� ��9;,�ސ#B��Q#��V��??���-֠dW������PLV��	^rv���q{2�������J�����nH]���$΄����c*w_y_j9@����w�pT�ֵF	��_-<bς��\#'>��O��7�s	��]�`k�
��紡Ǒ����o�<�y[�5#Kيo����xjeSkʂ{��Z�5[��F���vO>�����X�Dn�k�Wj��P�2+��e���`aj��*���*"�u_:�8Z�臦�6�bh��%�lF}tx!�������~�	�	q�A������jl�7y�m9}b��m�'G7m����\��'lO���K6���_��M�]7nc�8'�q8��>�\d�7rO���rK�rb��s�@�y�K)J�L�m�����ɨ6l�� )ax�ԟ)�!9R���Ӱ����Ge���hIn�*��Jd^��E>�v�;��N��m��vUf�X?Z*� �%ϲlQ��Wo�Z!X4�q�Sdf<�J�Ws���lx_Q�%����Ժ֡��c������<�=�����ż�\XH���Η��f�kة��z ���(��r9��#��	�������}���	x���͹����!�|��z�s���A��__Cm��_|�.:ݠ ��W"-K���'OI������X��DKR�� f�Nν��5��qH�}�V8�X�|�R�&�o~nr�1��$r�?�0�.ro�������)�׹"�}vQ�4.Y�ƹn��u����-E?�Pϻ&w�}6:�j�sߕ�PR[Ӊ�������v׃�����	�c`��*����`+B���=��N�.��W����檵�qn�B��U�@�ȿB�s��r-��(��G5�eۖ:\2��sF񆎰#�N�����M�i�,���a=�>^����^�#�␝�P}��1wO�j�	��^n�"J�M���g�P!Y��2J�xmW{e�2�Ǻ&CW$�&�
ͪn9i^L�~ڟ�y̔:e!��z:��ŕΪ?���H�,�C&c���dd��y�����6		��/�Pa�t�!��I���MK6��Mfz��lG�_��r���# ql��y�TJ���I����y�j�.�K�n���a6��9���ppu����(���\�pcˑ]9j��;���1�nYF�������U5�{`	v�-4��V�1ժ�$�#$�]��;��W�8E%��%Jgj�#���$��Z�uMa��X�D�&�4�6��A�.���,k��}z�z��$�~Ue�Kb���{��D
@0�d�?+#^{F�=y1��p����>_1�u�tf��`���
����Vk��|
 p�l�=�I�<��V�'f����T���u��?d�43��A(�XzT��[�R��E��3��[[���D�Y`�A�Į2U
���W��$�F)v��041�inf�¼�>�\���0i۲U뻖�'Җ���~:�-@���_�1�bj��V%ۨ�l�Ճ��*v8��(xY�PF���ǑjBE�4�!8q��̧`w���B
J
s��S���<C���/z,��z>v��+������t��N*�������6@�,~�y���C��o ������so�~�sFYbֻ=��L�7�Y� y�~�:˪��^@ �;��\�[FB<1�N?X �4���9@�w��	4h�H�;�0§vƷ���;E�����j�[����#`֤4��<(���Q_*xP4ê���b�)IH�������,@>:cc��_� �/xd����kUp�����e1�?B{>I(.���3htt��az�(��H��NY��¶Y-ҧ`��	S��Pc����w�v�Ȳ�!�릞F�7-J���Y܊�4�*��u�?�T�W|�g�D�u��=ۼ��>7b�I`��%�
���vu��_�婔I��L���q���N)��o�FK<�vK���FK��-{O{_�Ey����_'t��ӏ��C�˂�L��M��mfUF~�!��v��k(x�p�y0��xU���*TT�d��՗-�|��hV>8�������xr� ���&::��H��qp�Ӈt� qF}��6}'Iy�	�e\A����5퓤-`N2�:���ӷ*��"���H�Vhf�~�l랁�Ǒ��z�1~O|���VE�Vo&t]qA�������:�+\�!ڃ8�Px�<�1|HāP峸_���qh�+�9�`8��	�׀o��*  ��Q �Wj�8��'���ܐF��[�|��w���,}���<Ґ*�K�
���&g[��N����^�{���@��g�X��՚�2o(��������f��,4n�?F���ȱ_�K]5"�{��ݥ'�0�m��#쭃�Z��q��)���;��i���������{m8�y�w�ߏ�3s��}ｮ�>���ܥ�ԁ�S�k�6yW���.n% ���Ħr����n�SX�ð�?���A�~����Zsv��ߵ�خ��Q���еK#����X)�Bv̦��S����#N�Cv�)U���|>��������{i���B+�~�x�A�����h�}�=�L�r�9�Ŭ{A�8��b�|�;���;��{��j�v�ob>yx[9��N�`l{�0�����,�	�1����I�qu�P�)�~�XJ�"�g=��)V+�ih'�h��-��q�K�q���L{�C�[!��"�?u��
�O�cU�W��An�L1����w����M�W�G��	R"v<̂ v�ū`�I�!Cf�q�c�ZnE�i�	�}fg�Q���&���>���f4�Pwۑ����g��������L�Ǹ��W˛dK�$-ר�M�{�u7��7��UY�\ҿ1yW�]�ʹp�r�H��'�p�p�=�ܦ�܅���]k󾢬��C�����$�����ޥ�ݏށ#pQ�c,kQ�a3@F�v�5�o0Ͼ�8c}�X?*b
.҆��3��,�dM������'oFr���s]s�ovB��;����C`����T����c��J�~���{��B�oF�\�����H�)�z�<_�L�h�J]��[�|o�Q`�漮�A����e%+�Ѯ�~�=�B��. ( ��Y��,S��j�Wq�d=RR�^N�<!���g��ݍ��%��յ�t*8(���w�h��_J]�J]��9(3��c�;�����u�'A)�z�^�&c��o�71��t����hC��u]�:P0T���|�#oo��J
�MG��_Ӧ�'c��b�h�ˎ�Lhz{Y�d�ʇD����A[�Oܙ�e �j�y�o�^1�+���?oƾ���}5]/�!��-y���$�#+��	ՎIa�y�aC�"��&��E8s���p�\���+�<`-��$����V��)|��?�v���%V[o��|�y_��I*Sk�I�S��@��Z:�j\�uy"Xߢ�$V�+6�������?�9��Bk60��)�+S{������r@ٯ��M��/U��Kɑ@��q�_�	5���7����(7XL椁�����P}��z5�����ҭ��&�^��p��q���G&��$*L٣��G_��~($��q�����?�=��Ȳ����K����Á��cf:s��&-l^�d�x9Wcd�sV0�0��9�jU1���3�C�;���������
�g_�-���.[N���M�/Tq���J�8�E�3	��	�.m!'����i_�v�GA�d6��_�5'UW��
��x�"+r�r�v��۶'3�,�B������dH�V^m��&�M�������y%�6]�9�5������r؍��Tnm\�E��� �w�����)K�$�H/�0�Т՛��7�F�(��\����������uk�5��bj����Lj����P3D��+��뽓Y��?�N�X�r�p�E��y���c/�Gh�~�"�j1����%����<E�.b �0�.Oq%
M�ݶT����e��q&��P���6�v�Z�ok����uJ�2]�Zk(@�,~�nNk�Pn#���,r*�K��$��/�5L���ŗ��Mߠ��k��5�B�-�D�Bx5�����[�d����R�f�C��C��j</����.\�_�/�F�#;�I��mcp�g�� ��PIr�
����Ö�����n��J�G�9��m"8pz�l���t$�Z�KP�3q�_1q[_�wߝg��T�uj���D�W��'in5Ӷ��#Z]9t��X?7O+8k�=>0����ޢy���q��M3��R�(�����Fڟ�p��E�u�G
f�|'C��o��њ����I�O�����,d��#��H�\2_�A5g�n�\�EB0X/]�`p45k�:��*���
�:y�[���d�4���/��J'�ejʥ���@�.��,���%jk4���,�5gn&#�0��mO��5i7bbu���ޒN+$�`�UwG�+_l��p���l�e
�i�0�L�^�l�b���}���# >Mm�!����7�k� ����jG�I�:�B��!�+'k�0�]� ]ڳ~p4+�,`�,ݝ�5*<�y
+����U9S��=�hɷ���m����%��!Lv�h�9��mL��0tv�с�r��
5�w�Z�ݖl���^&C�Za�E��e�9:��2[-�oL��Uc=�MPQ�9N%�k3��"i����#a�{텞��3W(I�֨s�;�̘%
�I��_̥M��d���s�rרY��wJR�.�j�Q ֨�����^��/9X��'��U��X+3�y\�^�cw8����kλ1*�D��b4��g�����ǿ�q��R5�텂�㉬@�ω���`�	W��4p8y���Zm���U���lۇv8��
��R�ҞEk�ӻ����n�7z#<�W��Y����ܷ�TT.;#���6�qڵ�g��?�����G�G�T�6�r1�O�r�ۨ�4b1[�;�h����c���-���ښ�?�Z�
��E�tS/lh�15����� W.�a_s�$�b��f�+��C�h+�n���]%|7L~�<�����Qk�������\Z���5&I;-�&[�'"8�J�@D�����t|�.�����&�I�3�/l�V��a����3���W.>y-��Q��x���v�}Q'��x]�g���Ik���C}������;9����靶���m�G����픫!�
i�ۺ�՟�)���33{��i!n?Խ@'����2��@vd����{ڴ�1P@*���Fc_=��i�y�>r8vC�/}|T��^��0Q�`hl8�����;YfT�W���;8�/5bv�,��e!F��@ݛ|�R^����~��讍#ec�w���םg�>�����G-/?Y �4����@An��BVe&Yg�-�,�ܥp��s?���$��[��.�O8,^����W~���%ٟ[,�ȱ�HE.\St]��Qբ����Ft�o5��u���+#�C�������*�r�j���,�YHy
o�q\Ox�K�|��PoF�R�Þ���O���`���]�٩K���,��FK�0�Y86��-V`�]e���-fe��~��5��Sʨ0�o�Oj^[g�?�ɉ6�������.ZTiٛY�;�H�GY�F/~���I��'P���c]��k@X��z6#�H�F�򄂏|{f��~��%p�^Y����߂o�ޗ8���&Qڽo��ީ.�(v��J� `� ��^^�涢_��@5u�Ux@b���C8L8��_&�P��:��T%bj%�hw�%�x�N�h���<2��;�����y��Z�B[��:/�@�Б�.,V�arp/���XXT���Q��y��,�.ܥG@�i��\$d\���- �_��|�!�:]p��t��M6-;4w�+$��T�;����M�v8O$\d��������[B{׀!��8ʠ$�[�� �G�Q��4��x0��������l��h��q�q�*/����l���K��fc9܃P���
���U����w�m@!�BG��Z� �Gjh&�0<��x�+D�����d-+��r?&Znz�ݰpד^���`�o�M�Bw5��	=U�h��C�y��޺�ug��)�e_"��0�w:6�f�v=}v;0��1�1r�;,1���-�Vjj�_�O����}��-Α���/���1�=��߹�7 xpD/�?2Mb$�mB�� �[I�}q��LhC��wo�ͧ��^ޤ۶m���(�z��C{����
 �Piý�ta�ոX��G��;���8vv1��8

:���Jq�Z�Ѽ=z/i6��fj�6�2֦k��[��:�?4����x��v�����(1'�h�f�*�e��iZ��M�ct������U��A�+R��=g�6��7Os��b�tj?���)��$8-q�9����!�@�����'�0�R�F�w��}ۙ�%d4Dz�����\}-5'�)�}����~����f�c��j�-+��-�dk'��I@K݉�Oo����4*6�ޛL�Oɘ(�{N��V<uՈ���P�=֧�)��h�_֕��Dľ-��G�������xK�_P�/9r]kX�fl=vOԳ;c.���r5b���N� J�Ku3�⒰�\�fZ���U0Z3@��bj���_��D���;�1�.����A׼�������Gm��l8Y�,��P����7��=��^����&��h���pDƬOJȰ���g��yd�(N��(�^}����Ml�"!�<��`�����(�ؓE�NvJv�+��b_�M���#߬�*�u��}�QA�p��*X��n"U�������F�l�SZ��p�r[��T\�j=��ܮj�7U�,%�M���=����2'�o����5�����p,7�o�-zs���D��H�w�w�x�wE��jY����g�Qn-��D���NM�����v�t����]q����-
�+�p�̵��v����~ (����ő�ݨ�_b�	#��~���M5���R�n[��)
+E������������닖[�%Ih�,_��C;bI�'�%|c���a��X��[������~�5|EA���۶�]8:r��狫^	�d���t��մ�v̺��Q���m���;�R�hR�W�[��I�nJQ��H.��[^a.��/��DT|n��7�{��s*��ll�GJ�uX]��.��	��"����˔��Q�.d6HO���q�j�6� mq��]����B���2���P#x���g�6��p�T>H�����*̳��������(g\��-Σ!8@cǈ�� n�Ï��~��A�,���1b��q��:�I�,?(X/�Q�`���j9������<�>)\{cY7
�'�6O���"b y�C��2l�j������~�F�]eu�ӣbƶ�����fõ�OB���(l,l�k����%Gq|�-�IA�;��Lr��v=Wj5s����ڵ��c�"��آl�ԙ�v�[?�[��H�}��o��`^��,)񷽊��;�{�u֮(p���,���yT�[��Q���Qi���56�~B/6���#���	��A4��Y���ʆ�( ��iY*��7�ѫs��O(4*�����5����
����tݪ�a�������|��4^p?9���{ɢ{�FUvEC�"Q�RӀ�d�SaMf�yt�����I�|�̾��!�W -��TPi G�k5\l'\D�ͮ���]���ã�w���{I:�9s�G�[��s�u��9���*w�ת쁼�_���{�x��pO�Y�͡.D[ɬq���AS�Dt�I�.����ŵ-���8+���e�1Tl�=��Z�������:d@�'�ԙ�vC�iOhws�p{�Y�%�>�^�!TC�[��P:�3
�����+�iȃ��cF��R��.f�4�$#�<ԕ5D�a��w��|%L��y���GF���0��FZ�ѡ�ei��t�ms^v�Rn�|6C��g��<�p�Z��L��Q6Un4�\��������QA�9ӗJЀ�f�6P���:��Y���'�<փU�&bP��Fgo��x�#@K}�}M��H�q����V"����C�ڑ�������HI)1���թ&�nV8�������4 �JՐ�u���C&�n5�ŌbZ���!KG1��`���#�V}5�8����A"zM-��p���R��o��et?��j$̙Wl�Uz>8�?���2�.O}��[:z���>YI�~Wl�<���yAP�mnq��J׍�'���􏹕�k�d���d$��%�8C��h}��J#C�ы�<�0=��V�hQ�A�rC�ȯBp�偲�&��d�5�����%&���d��:�S�Z!�v۳2������Bj8*`]�9��WA|��t�	��m��c��ʥ�2�t�V8���Vl@����]���м�A(-l��YB}s�1Se@��[a#���xٯ>���j{M�n���%�gH��P,վA 4�&�.��+6'�A-􎤡�iť&�|j��j���_�Ҹ���}M���!V�V��Q�F��~I�򖕯N!h@Q9��m��B�%��	�`^wB\����v �m�C�ϒ��[��l̳���R��Ů��eq�e�C��+�WE|� yf@��#�1	o�dj����MM&s�Kl=�dM��;�����/?3$z�KC38SP/��ⲋ�����G�)ȳ�|X�6d��h�f\ �����`a�e���˘�{��������˕�5VlOBA�!i�k[��+"ޚ��%�C����}�4~�'��7�7�P�]^v�0hn��D�Ql�\ޢM����xV�����8x�"��(Ph�~q��XK��ҹt�j��0�a/�zb�����h.rԪ�A�j}�Bv���L�B�5������������6�> �M�������]��� ߬?���mcT�}�#�)��1���R W��	�~}��������\�^Q�%�%��м$ʿoHx}���W�J�%��+[���kۦ��tG'�݁�d�4�(�6���q|��LT��l.� �4#-���v���\Vc�_��漵���;J�ftɀ$az����Q.r�F�#�.,�/�h�p��?I͙V
�o�D������;�?��ֱY���G��\�.g
K9�U���ȉ�R�*H0#��\��ݞ�~W���q���v�JH۾j��o�E���}a�4���J]
����� .��|C�.^� ��2q��l��>Z������m�+b�B"���{�<�?�=�w?�G�1I�	��������y�(�&{��w�}������]�!�2���j7*�ڦ<���'���H;zA4拼z[][�A���Q��ݛ��22Hh��7��|?����,>�C�1��4gkJ'�\�=2�3�gBD\T������R��=&�m;⟻l�	�\�:��g�Gښ;�M�b��lI�bȾ28st�l\yl�I��N�R�Qض��k��<9���{n`��/-.���/�0�lq���t��&�A�͚ےLը��Qd#����yc �w���P�P�n9F��YLv�P�����ԽM�q���C��69������$ɩ�0���1�|Y��WK4�p\�[��L���T��LN�,�����{�?�ʕ�ъ�ԯ��J��6��I�^W�}$\�H9~"N����;�J�SG	�;p~��HOH�Ƨ����;Su�u���:����+$	�AD{���k���m{�������xT�k���4��d�j"�t$�˂���}��v�L]�u�Oc����F�'�.��	�;i*e+�)���a�!���
�?m^�u�v`l����U��TįD��7��M�H9Z��/�DR�G'�{��0�Nԯ$�臒�9<Voj��e0>�v>8}��	�5M2�A�ӏ�C��m��ӫl�ha�d嵰U�B�7����:�?��Ka�(����~2������6�V:n{HV�3�E�>V�ƀ�����?�9�_uIFf��5-3|r��������N�0M?���m7�\}y�˺i��HK�I9��y0��8�hc*k	2з����U�\�s�Y��q�&��y�<~�Y�J'���O��!���+G���n@?����
M��6��s'����L�QLa(N	���Ŗ}�q����C�R'"�l����ȯ����6���|_ܓ�\/�t�yS���iD�������(�on��I<5��Tѕ�\F��iN������K/�b<�R��l����8�O�9)"�bk3X  �;�ZQ	���q���Ћ/~�)Gk��{���3��Y���	;�m����6�?m ,%"�su���5�F�����݌ml^Ƀ���M�kng!�8��տ���˿� �ݔ༭�Q�j�:��&���<Xx{�)Z�9\C6��G��'�q����7��]���?i�� ؐ��Xo�y�z�����+pj�G���U��Rp|���'�$?z� {�Gr�Ә����8hǟ ��h��?���M0��kW��o�����z��b��rޤv�BXn>HB�j#��x=a�OF�@Ny^]9j�4��Q�Ɋv�>�;���0�2w%E�D�N��/W�|A���1RÒ;��镲��Y��
k���5���X	�y�q`�#���ɞSk��n�~D��NJ����/}�q(!�g�
o5/�l�Ϙl��/�����ݺ���e=r�r����{�.�Z���u��JlUX�g@K
�s��5��^��{4 Vǳh�ꃢ���+�_E+���0C?<v�3����
�Z��,�@�N�?tzZM���b��jB|?�OjM|�Y��)�r�7Û�0�)�C5ܤio*�889�%��Ց h9�?cf��Xx�Ze��[����g�5�6Q��������T�	7F��B�~�㡳1$~z��b�S��Թ��gz���I����ݎ�j�3���߇�} �F�.[�4��n�1k�ͅ�|O0�	Rt�6�X�M�-�f�~��g�^i��ƚ���O}^i����*�b�Tu�'#�c�
p�]z(~Cc��P,1֤�7��u�?F��Y>�1���&���)��l6a��6 s�����,"6���XxLB����ޤ0Ք�z�+���ɯ|��c��=ۥߎZ���>O/�A������� ���_i�n������S.� �-�E�Wߚx���#��$n����/�[�e.d���,P��.L�T����j�m�g٬ttgOhԉ��<Y���D������LL];�_:3)j�_S��ͷ��!�8�Tw}kJ��s��d�$3"������媛<l�ZD�zp�W�qN��t�W�s,~��};KC�"�M�Q��A���i7)z��	@5�mz֗R�Y��<��'$�Lg��/�[4�))�����=1\��r�4b��H��πft�2HE9:�	�, �
��f& #MyI�%�G(�25��h�|�|Hʜ����;qڷ���E\�̭/����$�������j�7p#d�1���I!�[���_�m�v��W��gp�fg?�=~^�0mv!3�1z�&�R���'g�.B�_�L�9~y�i����N¿kH���P����rG����յa�i5�F^vC�;5K�d��s]6;��7l���%Q)\�����ғЧZ�\��w�xH�"ЏJ��(�UjҪ����D�������*q;>T�#کD��w15P���:��C����/��~;�4G<��A��g� ~�n��+V�{'�M�8�5�u4�sQaỜ2�j���2�����Z����M�.u�������}߹����v��%<Aʒ�������պ�B$������G�{m1fJ���<�c�z�Z����|?	�ј�l��Wbe%h��`o�=C��	$M;���F��q�!��B����79�	�2ʍe�� "����r:O_�g
(�J��hͯ�4񥙘���l��n�}�!Ͳ�����0�/��Y�9^�P�(9N6���+RNm��)N��?��j����QF�����"��7K _B��kòt��Ϳ@ MT{�_sh�6���|��I�qp�O�mi�4O�PhȰ.�ڶ��G���x'��rY����È�In�
�}� �w����3�;p[P��~����|�0W����",l���T�D  %���C��.,���i�S'�/#?��b	�]�G�RyI@Y���åB�q���Az	\����1�f;\=����X0x�jrl8�r�b�pi&o��	�l�v��Z�_"a ��}'K�����8��9W��D`G���E�W�R=n�5
��0;�{��pv�-p�� ����~���t��FFl	f�n�rP��@���>Br�J�<�p�ټf�c�.�H8L�+E��:M}��Pl��f����0�m�ؕB6f	@�r�s/ �j�Up�f��n��vh�;<y �$�m��^����|�ur@ܧ&0�fe����wT�E�"�E����Z��4P��	׌%%Vet>"��XS�ĺ��u:�޹��h+���c����W}�^쾥U���ō*Wz�KW(�:\j�/�(x=����r���פ>#���^�*D$3n�wϖ۾������Љ����ǟ8H_$��k�-M���~�{9�)��!��nno�k+�,�{�W>��ge�]ʵ�X���m�I����{���H�46�z���2:A�q�S��g�jE����GkCu)��K���4�J�}�Å�6fb�(7.�E*�IQG�:�`��O�}�s	���=�g'�с.AC5{N�><X��F5�`6��UHOH+i7!��,�tK���Z�a��SU��0�8]sIn��S��0����u6��"�
��@��j|[�����	��V\�~�C��5!Њ��M�penZ�Qm[|����g�K�^�q_^7�K,�"�3Sn�a�_��e/��']%,CH�F#=[!ϰv��<�k���hYYX
��a(�[���z�F��ATnR��|,LJ�>z��Ց@��m~��Te��T�K#�lm�:޲�Q�Տ[��?�VUf�F����h�Lv,،L%�E�p沑T�PھlKJ�􏽺α��d�����7~)�|Q�s�3
=m݃-rƧB%�!���W��js���u"|5`�ٛ�*R;aH�mf�5�g[[h+�Wk�q�[�Ӄ����?�2����얦b����]�a�3��*!{
�e�fxZ���-��O��bi)�A�|�7�b&8/ȳ�0����9O6(#���=�d��z��*��{�Zz��W8�+���)����?ߊ� ���^Z"��l�7���{˥j �W�?���"��,�0�JK��:�����MI��=�$�R�\�`����֖� #y�.�"qڮ0�E��+�>u"jG�ׄ�����8,�K�wAq�W���}��(�35��`��v,/>f����}J���U��	c�bF9:E�@�eC��o�*�B�]�H��ԑ��ɹ�@#c��	��jR����i��䘭��O+��MW���MUwT�~X����m���/�6�wk�/���I���@����a����*Aƺ��;��l�� B�� �c[[Žs}Yz��Ҿס��l(��R�T���Luj�+�!m�ͫX��7G;�6x���(pu��u����`Vw� ٪|g����ܿ,��I�����qy%��c�#���6\v�s�lX���46��%�o�B��%��_���E#-��~���RŅ,��K��:�@L3`��dƉy`��q�䴁,�y��+qnF�vvs;��֩�f�ힽ�t�j�n�3���"氰�n*Qj��1�)�Ѽ$9��]D(ӆ�d]au��̓����E�Z��o�Cd����C�mHxmUT���ya�k���Ʌ�A�\^@�u�U��71wnF)�+���!�`KRuCe�Du5`0|��!�[�����K :x�P�Pś��ޠ�[UU��1�Q��+Ղ\4Z��A���+)�RY��E�{2 ��#r����!��"m����~���$!:y�B�$7���d+��v�P��=?���&��F���	1���[��+�ڲ��eb�_�H�@�^ �[wf���Տ (Ud?��ũMkJAa����D��\"�6^� ��' �]�1�ؼ��oOޤ��GU�+tS>*:DĻީ�^�!�n�-o�;9"�
|����J���Wg4ԥ*b��UP��#�"�j�{�*�{jn�6�4c��"ԫ��r�����Xz㈄fw�Z��Fv��0*Èf��j�,/��Cc<�|��t���;U�$S�2�� �a���f���(��k_A�~�\�a����!J83 g�7��`�Oj�;8��f�f	9�g4�-0�nXӓ?�;�5���ܵ�=������c��L���[��K�M eW%�����> �o��s>8���Mp1K���Q+,�����/=e`Q��G������G��U�ZOv���^2s��qU�Cx�>hψ:6DabT��4"�����M�D�T�\S�ׄ�{�_w�u��f~�~��0�/�U�=)�Ɵ`���wxI8DȦ��B=�������@�����E��h_�$W�B��=>�s�zYs��$?UJ�b�M��5� �[�f�O޶WF���+Eh⅀,���e��3@��4�v5��v���pkmi�^fXZ�V�!�,D�������W���a�w2������V)��b�>�C�>=;HQ��ݓ���GH���S�5,�1������>	�����w�T�tP�
��a4m��|ݾ�up*6�
��=]���{�JQ��dK� ������I����h"1"P�+��ƛϗf8ƾ-� 呁Q m�/#�X�7yo�� �k��V�J\8��I$�8�o��x_%$��Ou�������j�c8�&s}@�گ��Gr�
\��1{�S�ґ�-aF��kK.F%���BC�n��vb����u�w~c�hmw �T��4�g:��7ȳѯ(�v&�^� o*�jsT�@���m��{�m��H�O�)5��?b)��Z`-����y����ں=2�v�E����Y|�@��4�W�r�	/Ԍ��>$�Z�'#�R��!��yDq����=/1�F��F��9��=`�܌�N@����'U�`�a�NL��Q�Q���Ⱦ&X��E��C�Z1\�����;�W9�t~�\��W�����1������t��7���G~<��
�+,�}�/����B5"V�܆�'�S����n���?���b�2n�K���	AI��ӊ�Q��=2�=��g�'.�7m
���x!Xnsm|R���9��=��ՙ�կa�����J�uW~n�Pm/ ^��J2�����[_ƃ���'�R޴�#�XJd�kr1��$�5i�͟���1�q8��%��>B�NQ�������O��"��g�x��y��!4@[�e�!VmpQ ��	����v��$�����)1\�he/0�������[�Դ_R���z��E�:��ݛƗ�����ib�PLƦ�`�\�i��q8�=f*M2�,�H�G�k�+��)O��
Լ�o���%N÷�q���!Ny�۵���xx�~�
�(/��>�����zR��`�V���J���)V����E��)L�	'c��`:�l�8���dE���9LbDo�S�2	���y����~yd���X��i��w�.ϱ;��=D!}l���<�Xх��w݌M�����gm�lI)�$�||�&�x���L̪�����!FBΩ^��z�`\e��LJG�J�pAˏ��j�f���?
d~ý��D
nf�,�T �_^�3�!B�uҺo�c�X���PÅ�hc \b��$�����ϒ.��S���.�oU����D�Pr"��n��^��'�y���`4m�ιzI����l���D�s*%��x���=M%Ǳz)�{7��4���2���ᬖH�>�5L.�7��s֍�:�fS�	:<�3�`o�����Y�Zk��ՅD�����ɚ[P�RhI>���\�?�h��cGI������~�t=Йh]�� ���i�W���Z3��.����*���Ώ��^���4���z��\8�q�q?���9庀�)�y0�z6�[ۄW���>J,�������Sl�2OF��I�3��w����v�T��O_ц�G��uA��bE�
�*(�n�K�7 �Q�&��\}���mޅ:i(GKUN��6��.[C�|���`JYD�L7cK��$��yb������6��=ndo�PX;#���V?x!�� ��]^{"Xr��B|�������K{�
�?���V��IrЉ<?��������~���'.�-�%/��*X켷�k�Ĭ��";_�{���{;}C��.^�[Y����4����m]
?�nI	��*L�����	(ٷ�xOσO��ML�H��`�=�(�F�{��K�S�q�y��Q�V�a�&���oҨπEq�(���h�"��[K&�
�}�*�_`�f��(�o�w%dɒ�*؊ $���g��JDʩ;?�TD"�9qq���Ɍ��g��_π ���M>8x����X�փ���?L�Z���7Q&XR�8H��h�\���9��a7��",�4��rq���������t.w����ݓ���"!���09j%>2Z��i��B��f��V�>HЙ����|t���<�}���CZ�|]>�4�wga.XB��5��冲?ʘ�\~�S.[��GD�p
h��"��?9�&�E>0\����C��,��
}���b�:��Pt��=���}�Z��/q��v(��G�ǲ�Q?���B�7P�L��Y%��}O��7����� �qvetA��^
T/����1�0M}���n�Z�:]&pu��?$��9�ﶲ�m�Ah�\�W�Q���&���h��Rݴ��\�Rn�G�&�d�q��7�	�þc��&x�7W݁����\�.��L�55����;x���J�@��1	����s�;(� �e��-���ڨ����)�C��gz8=����|��e����aÅ���M\�C�sҒ��:?��8VI��< ��}�I��,HH�F���x�kW�9dB��ަB�	���>:~�Ok=�)	
����\��^YG~�ǋ�'yʊ>U�d�������р�3l�/K:�S�کŹ�X��R�o@�XO��9'�o��]|�G:l|�5�"�R��  �q�ATTō�G2ѝ��-cC��D5��1�/�gz�Z@܋?�@>� ��w8��F�)�������N�*�L+&�4�*���/�g���#f���˸4h�m,���9ѯ������]�73�ett��Ӌ��?��osfA��p�{�':��J3ْܛR�a����]���,�Ze��������<��W�H40�g>��b��'K����_�-�;�!򕖦��/m�\Qb����5��_	͟M$��%\X���]�H�J��VU(�M�x�f�	c��+W>��o<�?��U��f�ҕD�ѳ9V���9�Q�p�l��`l��M�,(�Єɬ(ޣ�{#�<ó�������sfF%ڡ��i������Vcf~���?�3����$&ϴ`@0H�$�Y�s���J��1˒�YR���c꒖�c��{w9�����*i���tj#��d�{��x�(9Fh��u�����7O���q0`�w�$����c�����7�*P�j!�']8��#�p[�:R9վ±v[�?mG��#j�OL{�����<t�"��2}T���#�*.N��bbe�����(�UΟ"/3�����?�~����z8N���%��{��
�&R��f�����J�\�+����X&)3�
m�ނ����cXDT��+�Y*83;���0e�e0���I��T�	/gR=^Ȧ٧\��ӧ��Ŝ	t�n��FL�L�G�q��#Y�ӃhI��8��iΪ^=�GZ���4�4�8+����ZD���*�S�r�!h�1B���\ʇ��s�~�F�rz F�<F�P�o�� <������^Xo�~T���[Il��A��2<���8`צp\W�&UWB=��V�}�]<;�Ŀ9j�M��آ���d*��c�m�w�i����z6P\N=�$� x�w�yx�uj 9�Ѵ9Z�!�H��;���76a��=�:�>�!}�Y|��6�]�@Q����_;]����٨���R@�9 ��.% Y�z���4��g��0��0���U�z&�",-�b���#ˈ}k"D�����B"	�����?iU��7�mO�I�&�G���*���$u�FF(������2C����+`ȇjhK���_�>��b(pB�+�ܧqY�i,����r2��@c%�T���>��i�j6�&��p��=�9�:~l�/%���o ��s���M�C�PZ.�{<�c��qI^h�I���q�>,3��īN�~x�A���W�`���%�Lŀ�8W���7ly��x ;���3��%��
[�s�����̊���7F�E��2/�דmJfF��`����R��ڐ��M%����+�Z�����E5Q���p�,P
$^o���1���[�m�h�Tc�F�^p̂����=d9�-��^�ܬ2�~�,$��=I,POH؟��%�3����
؆ʰ0 �:����\�ܩ��L�/HI(��[u��K�к� -�̗|I�^����P��l�BM�=/c�� ,���S��R%e��&6plY6x��yq���ixD�A�?�y���O�y��Y�O	��y8�̱�5���Grq�H�$�9y�NS�0
V��s>oc2�N����<�
�,��߲ᓚ��C�1��r�3b_nsk��f�P$i����M�s�b-����iW}����{�7*��1J�J����x���T��g`��v�ӊ�+��e���[M�J"z�WU
�R^O���CF�y.�v���k�oSJ.��p��a��3֧�L)y�tz�+��x���-�X�]ދI
�Q�,���5~�o��hs�Lx�%�_����#�Rn$)��-��b���//�A	8��5��_o�Ts�DF�`v{��(�%&����jΗ�p�.?��d�ݛ�J6��7/�� �sO����3�]\�����Pʮ��֋����]:_mX�F�fR�ҏ- ��$�Ѡ�5<{�k�=�r��}�E\��iT��e����si:Q2��
Z�4�Q��#���m� ׯ����j���|�	t����Zh���|����.6�*F�wl^'�,@�<=}�t��O{MN�M׵R�Lt���I'��2gq�K���o�T�Jz��_�}��7a^�P�-%��*C��,|l��x�0
F%6Jzt\ӿ8YB����u/x���>!��Ni�g�lj'x
�HV����iV������4�֒�j,���El�Z'b4"����<�� ,N7B�L��}��� #Eۅ�zA+��΋�,k.����&,�Nt;I�s��g�4���9Ԩ_ǝ/
���-A\��G}rٕ~��d���2o�����:�X����y�H��V1�`�6���D����yq	��E�:NH�1ǈa��M��Ϙ.Qq�G:��S���9 ����X�[���t5?}�����PmˉO��6k^o��_7�9Es��0G���>+�T���	@6����༑�$��a*��_��|�C�{��P�-Y���`������c�G\�foJp�����6#RR��[:��_շ�?��X�H) JJ �%1�tw׈�H7()�tΠH#�3� C�o｟�Ϗ�9��qf���z��������r�t`Z��$!���d�y�_�&�������3�=Pb*0�hq�5����2�u�v�z>7?KuM7������Y��7$���\�F�?��w��B��׽f��d�I�FL�'�(����o���yf݃� �I3-8��ټ��������p�7_V"e���
-y���-/��W_!>� I������ŭE���n����Ʀ�Ɨ��^vn��w~�$�PI'�a�1E���V����
�)�W���I�L��}%Kd�߬�2'K�ஷ����{�L �b)����%�(�I@���OnO6�t&},���}�*ŀ)0�&je�Pt�V���}SI����N�W����aS��G�ƫ/�&6i0�,8��O���GR���I
�O���6�f��2��x��b�I:枨�S f��`G�U�N�Qt�:O�6��3wh'(v��
-(�J������ڦ��!����7�g�u�Gn�{���91�]����s/BzuJf�u0��8�M�J�X���4�51�h.���Y]�����x���鮉�YȐ@ib����t�ף����u��"u��Ǥ�t�u��u]�,"Y��\I^�����M�R�7���M`RӰ�;�D��Ǝ#�0#���|e���e||�Xq ,ff~��<#Sس�J;�b�%���puq�I��*��L�+�R�&���c�����6/_r\����f���.���Nd�� �G�)��]�����EG�&���s`; ��T�̂���.���J��!Н��[��޼|��7�`InU��|J˙��x��٤f<�:E�ѭ�j��Y��M�mr�Q�р���Ԉ$����B���?4}��Ğƕ��;;�(Vcg6��r��Ӿ?�.�^�,�>��M6,i�� ��e�Vt��;��yf[M���?R{G�%3�<I#)E+['���h�ֳ�RG?`!�P����vط��A�t�������mƶ"LBL�dI����!�@�\2���"�Y
�[���)S�z��[��.�Ǧٛ^��Հj##�h�2�����t+���-��7L�fd�#-��������&�L�Y�:~���Y���e�(�x7��5���"��Z,��4��EwCͭ���/&�*@�*��/<A.o`���5�H�uL�f������2�q��J)mL/[�◐[fhdӞ�'"2����a�顶�������8ҧ�#_�� .���o�l=�����?�<�E���M�̵O�2x��"�����"����{�/y��l�փ�T�[](#7P�w� dA^�G�Vǳ����/�{�#�(,%����	�����8� E�ε��E2*�EJ��?��,U���w@-H�_������`y�њŎ�fR]�0>_i�z7���V5V�amLi�.E]�2�OCk2�����7�}�_�(�/��`�U���AS�H%�9���k �Y����YY�oG�GЈ��a���?��w�#�E�s��%>ly�ʘ�Uu��67o���tj�4j�f(e��I�/~�[9j����Λ�.�X��Cg���RN����gx��m�o�d����|�\侰��Kg]F"�Q��i�"CO@TKћ�jӐ��������e�����(�-K~�R�Ϟ�2w�"�Wә�(��Xy&�~�E-�-<�}��ʟ���?ON`D;����<�j<+���y��Բ>��1ʨt���=B�)w6DL~�4c�ʂ�M��(W[b�%O��H���F
!�t>��s����,����}�9+��أ������xs��=���b�*�VnÇ5?�K��t�V{������Htn�h�>���V�=��zȞ��g$N�I�M��y�z�i{�sW��ނ�,ޣ�t��R�u�_���8K9oe9t<wt�>H�v��$�ƻXUѴE�K����(K G!�|������Fu�>���֋Ga��;~`�����=��}�*��F=��u����QٚU뀼��zɬ��-�ׇ�Y��<��UD��S�@m�R�FC�������4iL�M�1vz�ع%�PN��o3X�������})���Tc�5�zK�Z�2�{��1N��>I^��v8�8�(e*�NL��c�@VW�����	����I�
D�9`j��뺬$_�g�,�RɨݼX?���j� ��W;��}� ��iY��U����p� d1�$���>�a�	 ��@}]G�1>�ڄ����]~*B����ms���k������G~�[4R*P��	׾�� ������sŶ�ʘk�М��������7RuR��D�)�asayX����n��4�er�^�����ۢW��~ś�2�����t-�v?�����hƤw���X�|�T�<p?�G��������ϋH��'�gQ4�:Hx���g��z��DfSW�K���?��K�B2^Z���J��X�^^���p�����%��f|J�0m�e7qo`�\��w����_�r~@mL|�hv1�X��0y �֘-�Z�B��L����h�7����,��AV���
'c��U|Pejq�>)��G����-�X-5F��jG�Q�uh
��ڃ
�HnE�w���,K;�fp�oN�zz�:�-/��Y�k\n�'9�
 J~@.�n�ê�y��谰x����S�̐��y��:'�,���5Ο���(4Լ^G��|F�^G[G�8I��UHs���o�oK�~:DQV���FM����#���F �x���[h&��]�9����߂�^�����8��\�=������	2$�x���:��4�k�,��f!⁉�!y{�X�揋_�[� M�ti散��h^y���B�$|w���V'��pӫ�w�s��ywN�й�*�SkR�l��\�P"4�Ov}��jȔӮX�}��T�r�\�����SY,Q$���Pk�[��:���T��5�f ���|F3�]��"�,�H[�N�O=Tg�n���!���[}��f{��艔J��T���^����5��?���^I���8����#*:�A5ج.:�M�t��v�.����ݽ�~�"�G�w�NȕW�5��0���p�U�־Ky�}�c���ư/3&/s������͗W�Ʋdl�Y�L�:��}�������%�q�H��nR.�:�wc�,~׏S9��ߍ�ϳw]�GZ�Sp'Yy���'�|"���=$+���z�?s�J��	��yo:^�|��l3�v*`���P�I�K��&]\V/��T�����e�`[��ԭ�,b�^��r	�����0h�y6F���\�~F,�#j�I-S�MkW<^(�4����Aē\'M��������
��z�3�B�Ii��q��/5�L|��*u*=�8B@i����teՔ��[��җ��2�x�.���\�|@����e~e10^B�3I�����7���{���������ׯW�f[���*uZꢄz��������ᰉ)N�3,��#���(�Gc�*
1�v)����n��j�1��8O�����ܯ}��O��!��؇��&�����}���}Z���܋�i�G��$>�;��K� ���d�B�����I�eY$7�#���9�xS�[�g���֐f�k;�MS�h)��M�J�m3=���}N`��P<� (�����5���_�
Γ���ꓪZ�5����k�OIpY)��7D�fِ���e��%"�E���l(�_pww����v��6j��uϋ�1f�`��?N3>�^72E����h5;��Z�f7�'q�u��H}�	��I��IW�x�Z�B�ў3*��GC����f$o��e$zG1�56��%��:�����iL��WYѦ���A���Vm�8��[�O\ծ�dq���;,0�Ǩ�k��,ö��ʙ��áIʧ���%�3� :�A��G��=1V���ׯ�R��ς9V�	���|ۓOԦ,0�r�+�j�lk0h*�����F�ܽ�SB_[�t���k(����L�}��Sh��3����DxA���s˹�hV�LI�4����˖���Y&��uϒT��Y�}J�Ϸo�a�������=�*���#�O0�gG��5@����{O��~�O�md^+*����yH�TS�T�b[5�����/J�m��3Ub��q�`j��M;�7u����x����X���2�a���9�����c���	�͇����{$x�ސ�	�H�D,i����2����Ǿ<9�GZ׏���,����'���<����w�~� �7��	�/��
j7?����HN2�(��?��ʉ@
�H_Yr0���&�_9�d�K��TI3��fc�k�~<���f]WFp�=��[���բ}j��ZOP��i�M�v�z�k�՛�/kv�x_�HH�L� h���?hw����
���oln��АrOݣ�'�Th�E\�/cf4�T�A�j�
,�@4����+��R�n��6Ɍ<���}//��(�iOҍ`?�_9�ă`�Ǧ�Y/A�c�7�j%�,�	���uw���py��	S�Kz��cۇ�t͍�`�O��h�c�b�t7SQf��[~IB��;���	�{*W�*`V����OZ̍�6tA�O���<�C�]�=�R��Ӹ���}���8���d�O5ĉJ$YBБ�"�~��$���g_vݬ�j3��I��O���	ރ&x᭖��c�F��đ\7w��\�}p	�ޡ_���PJ��]b�<���U���0��OҰLWL����DdZ��R9��8e��j��+!ƑUO�ln�m�H��6�q+�H.3��1�����Y߉�4���i�Cct����s:v_������2��%�X�y{�����x�0N�_�=P�g{�s��T�݆��m��?���tJy�"�v�U_�+���fG
Xn'��@K^6~��QՎK�ҝU����Y�z-�e�/���%�L����g�WU�d�xsդ!���+ǫӣr�䤌���n�������v+��?�ug�&��eKʓQ&�a I���q�@��M�}<��D���}j}8�ilb�.��L�����]�ׇ����u�^b`�
���'���G�,���j��g���?|���ﶦ�����	��<J ~�q��d7��Jv��
��踿}Jh��\$�������Yc�MH�^��%$g\�QL�Q�z�gT�|���j����ࢦ�Y�����	v�m@�M7MC#��x�;-<�q
���]U/��!S�y�����V�m� ���C�Nxa
G������J�/�|1�^���2m�c�g�|��f�iV�ލ����&��^��2��{�c���d�@��D� =?�[��,A����`�iz��eAǂ�5���󼱟����qw��J�K圄����Ր�{g\M~��<�Kٷ�X�����q�~���y��n�G��F��w_�ee%e����a��l�Y���a%us�nh�ޙ�ܕ1�+'/%��%�ٞB������|��vS?��&n3����+�}P�$;���qCGx������5�/}������A�S����]Q!J��F����X�8���EeC$qf���=��= �pV+��"U��kKs�ʜå�%LH��(~��M��Rw�|��7����^�}}j6L���:&��K�� C)>� 2�+Dq��gj V��C����h��������K�������&FE��:����:t|:7���r�;��s��8��Z7��F�����	\�#���u/VR�g/�?U�'�J�(���>tL3��9!� y���29�	K�Mi����]�����Q�O�����?y���)m��^(��Ћ T'��W"~���f\��y$��++ �@t5���
�h�-�.8꾳h�gA��	!ΌW5��%�\����r�b2c)J�i���t�w���MH���R4~b(i��~�7��W���{��Q�-,��Qx�W�}|887��L��#��E�w���q@`0>)J���V���K��nJ?<���x�Åu�0����N _O�YX�y�ۗ��_�}��, Q��m�������a�3�Ӄ�'_�>�o�����?�
��R���ZC��*��o��z�#�O�)��^J�Xrb�t�UO���rk-N��m�H�-KM�_٭PAm�p݁J�''�	c%$�y=|�Vc~��<��%�)1(L���7���fe7�){���>�-���ԛV�<�� ��%���'�0��ZD8�D{ ~ �|I�u��$�t�o���J���Bw7Ý��2����f\�ᙼDݙo����jw �B��:ǽL�f{�>�Y��l��s��nsO�}k[q��;J��M�}���bS2��)y��8)�R+��j��$�M��-(e�*C�auo;�ڔ\u�A�Gyx�Ѕ����'��2����t�����j�fd0�1eg_�z�>V�u0iKs�/S��+�������7��{��� ��Wns=Ɏj~X��z�D�v��������~/��J���m�i�q0�'���[�л38�Wz�5�^��gH� �J=t���n4�k�0�x��%�F�m�@P��[������Ps�"�Ʉ!tR`cʭ���,N��Y��P)5�-fz�������9��JV��4�}&%�Ɂ�T3��TXt ri��=�m �3�H�&�iI~�d����ή^��7=;t�$�Od��Q��]�w5G���'���D�
}|<��R5釥-Y�N�@k9��}�������M�/��n���cr��c�a��nx��o%yT�n:��Ά�E���9�'������-	7p������U;�>x�C�A%)��9|�����W73�u��s {����7�/���|���`�y�h֫|Ļ��}�W�����K}x���?>g���H�lK/���~A�5^Q�@�g���֧�a�ۀ���]0
hh6%��K-�8��V�50�(9�o�ύ�ƍ�׆	֌ȏ�a>ly�%�x��Š���A�''#蕎.��`�$��U-�Z�Oއ9�~t��%�J����I�5'�u�טVQg��5~����q}_ZJjk��;����
��mg}���	�J�W��i��C�С�����@������)6�a4p~twfs�.���^��������?���5�4�D\o:p��^a@k^�$U7��C�%�qv�
�V[+�1�n��뻩[���n1��~�y�{��gnvn]���6D!w�_����u��k�1�����˪07(�MҳJ�Qh�u��;���H0)�?jq���/��a8��k�&����C��zFD<3W,���ij�}ei���w�e�?ӧ�br�w4t/�DU��L��q��U�#mGD���Y	�����j��[�N0�h��Wb}��t|�
�|�Ed�V(�}�Vy�K�/y�V��J��R#�%g�R��Y����l.���y�.Ǚ��Xк�v=Z���0P� ������e�6f'��&{����������Ex��џ_Պ�O�'P��2��؞`�x�M9A�lv��c�~Ȑ��|�V��7-��z�E��-"V�pD��Z��~�cܔi�/�h2�$݋[H1-�{�bQm� va�B!|ģ����/�4�E��*��
�2s�%<i��f�����|6ͷea�_O����F�4\��3�ȒKN�Hص�e2K�����1%is��5xv@-��~��`oŹ&��d�%S�;451�S���X���`
SR���9�M���H�J%7��]�i�IT��f.+�E8�w��2��R�L�_�\�{ �}���{i��_�VP��z��pFw�Z�Jr�������4�,Qm4��GD�F��z��2i(�UK?�,S\���!6��FT�M���ߒ�};���CD5H0�_-�&� ��O��buy���G�D�{��K|&|��lBgl�Em���
?�Wdp�&��Ѷ�"���Y��f����ֆM=���z�����i	i�8.�G��G,���rij[��m1�ΝgMU'�|.�y�����;fk,���_�Y���	�M%C����2��uP����C� �<<O3��p���΅��p򀫨�"�&��m5���D��#�g& \N�,[v�uI�zA��5�����"G���W�����ؠ��h�K�G
���+����qi����~..H%��=���X���d�|�W��=�5�(Ӆ�3ҭr%t�.���s�Ua�5]}�mY,9f=7z]0S]R�R��@����?�m�W"�vG��u�l"�N��8�S����m[��<|M���W��E��(yn��
7W֥D8��I�NI��+��|�v���<�}�����?��f�_b
�����Cn+����ݹD��nz�v��	/U1��V?��U�A���4l�砓R-�R�s�q?yb��>���.���� s[w�=�Ӻړ]\�̀�x1�_x���l'㾴L�`o��.�G#�j�����@�o����8�W��c9����u�N�l$F�7I�Y��O���s=�����1�Ewv��܆mшa����\���pT�z�wh�R���K��TU�$Lv�<)�k�Q�,!}\��h԰���Q�0�~J%-��'7�É��`q�ΛL�'Vދ�%:��RA�@`�6��Ҩ�\�d�*Y��}z7����ZM����A6�o[7�v��ض���jGJ���Kk�6��T6QTF��ݯ��L��#璘�V����Y�dԕGo���{�y8�K�'����i���!���~����^�|b���v\ǵ�����K��`bnU#�/�pBԾj�Od�$�ٿ|ǥ'��>)���]���x5��m�Y�\9#�ױ�rr2�l�����Q��ш�A��B���f}m���q�
M�Zɚo ����#�Oz'��d���t��
������;-�͝
���ZЀ��/�K���C�m�,��|�L
�P+m��2���ۯ/Zn���A;.�{>z`�\�ED��w;�'���KV��E��a8D�����g��R�Έ�ň�޷��n�2\}�г�r������b=xw����t1���O&�+���dn������~����NF�+���K좇��Q�_�舿%ELGZ�n3B�zn�o�dD�/�9�,7�A�#6��
�-:J�����^.���=�^.nr���Tr"~:s̛�8��	X6.﮺�Jp֑M������V�t�8OT����=��9������n[I�����ͣ~[��#�x�~��b�E��Q�,�p�0�7\��������C	���<?1�=��)�[���!��U�z9X��
�����S�`�Uj�2��h�`�V��OJT�$b��������8^���{B�Ube�h��rgP�$��$�Rd�����lԕ�^Q77���"�݅���e��I)[١�띔!�g)��_���!�������}�]J�lm�S�8��(��*�E�N�A�^��~o�,����{��f�
�<�� ��z��w��/��/T���`{j��Q\o�+q���6Hb޳��S9�[:����.\c|���&���3\�[)9�qE���q+�!�\4j����ܰ��C�Y�V���y��Q�k�
µ�F���:܇�Ӡ�:����s�$}��'�Z��({x]�M<w��7�h�H"=`���^6��ϩufɓ�Ӡ�'�+��+���7���li{�)'g2�=S����Ц,�z����x��;]���%�& ��ȩ�dp�2�Q:����{�&	�x�Xh\��KG�M���3���j�=������-B���׃�����=��7�m�g�w���O�fi���d"���WAc$S=��|ֲ32�G�
�]M�m���~hp/h+�M�{V���a|]�C�qZF�tWh~#ݗ%�8c��Z>�m����<����:��]>�pz��R�z>�|�������]?�܈. >�!A��r2д�Ho�
1Sד���a�S�����>��X<�QJ��I����_�������-ԫa�q�w]S�����{�!� a�h�9tq�W��bǍNӜEa�ت�&w��k���$;�lW�8�1oG��_=��ߕ��o���Ii
?k��� r�
���~Xn�����J�}�J9��.����
F�M6�����>�8=9�sF�W�3��c���K��֐�K[�v�l"�p;�N����M�9E�(�z��A���QО��� ��u��bF5�%B��X�)�~�`���:`�U��X�4wg�O��zϧ�s�9fu��&\��;S����av9I�#�'����#������.�����;q�x|���p�6�s=�o�bS1�G����Ʊ�ZN7mNGG��(��G��헌l͵XW�r�j�v������hv�	���*� 
ڠK��HɹB�c��c�sQ��cT^}2L�k~��|L���,��Us:�a�Ț"C,~��J�<�f��}/�k�i5=�v�9]̀/{�i�w�ϗ��	�@����� K^Y�c������'�/�9���6�R���L*��[y��.���P_�n���sп�&��oq�]o��׺u�s��\?������7p��R�V�\��}����+J�-ɚ6eL簋�B�Lz�x�i�{瓺Ք̝q�r�䛛�	kRN�Wp��_5�c�_���aV���b� %�Kqu�u�J�Ю��_�1W��Q�n��9��.zs��'��
��P*%q�������J�G��P�*r��n����L��S�^No���Ы���@��W�g�4�Y�c׾��T�y����	� ��w���U'%j9��D��+|�7EF��h=�+F��lLI#��(���e9vhחϭ(]Eآ���k���b*	S���T��e�C��ޟ&C���j K���O��(A�bP1�����2���U��=�"r���^o��-�Ih����P?�.��U*��F�H����bF2t]�#�6�� :S�Iu+���s,v��8by�9��
CT�B�E��Q�����t��;s���@�� ����d�!8lg��=}�J��s2j@��q�n�Q�kQ�^�֎8��m���(�������a��SWF�Uk=��f��u��%���3��+��kY��H$��i���g����g���5	ob֫p��l�Hv�w�^�ބ�����3�$ǆ338�&��򆽯`[�Kg�,<��E��8�^;^i7I���Y�}�Ӹb}i���JRT���@U�����қ�R�3SQ��Vo�+��y��:��	��]�s%G�KF3��Vj�ס��o<l�hl�'��l?�d�(	%�Qds����-�|BI�=ƈ;�E$䶃���O���z�D�,y��Э.$���~o����5�����{�����J��"�������LRꮁ���;_U��*Ŷ���j�{پz�.�
���M� _F�����2�����u2����ꐎN3	���A��jf�7�e^�CH����Z��B�
Ɇ�Y�N9N�7[����3�w�X��w��D���)]�>з��KLxLg��V���=��dhByC�P7�P\�\���ۜ���=��p�݈2(�������*!n��ˉ3��t�C^M�;zvB(M��u�J!�2�(���
/�$P�L��v�L���햺���}�׈VAN=;'RLa3�5�7�D�,�p�W�{�h''l�,����`\\��${C�I�,uQכE�������c�1����bb[��Kk��5��I) �xD��{�'�6����"=̔,���e%�?rm�������5�"d��i��}J�@aaҭg`_�S�<�diku���xz\�Ѥ��eP2vc/_~%G��f�L��W��>m&<d!���󡥖�!��-�g��Oc���c�K��1�|.�(�D��Vz�9��
�廦�q��P`�~F |t�%Z�_����V��ϻ�?��0[C0%~��E�X�Z���O������P��!�?Ҳ-�[�����\|k��2��p��)�D������cn�~r*�"��&�@~��㾯߫��ɬ�I�K��e��_�C���|x.�:�v�,�?[7�>^�Ĉ�R�K���D�+��2%��d��^�:��DRy�"
�|P}���%�����-�bn��Z���@�`�](�M���p(��_�й;�t��C,���k�O�����$�X�_2inE��	{��Wv�1�ol�~�RxN-Z��D��%k�9�o�`{u7����w���Q	l(���m��j�z|'X��b���� �E�Ho�(9���:�e�O�CIZ��̏Ԯ(��c��{e�1�����~�2��rR���,k��X@՚���ǁ7��2l�1�O��Z������8� ��r��2����Se���B���4M狭���|)i��U�H]r�/ ȯ'����̫���?�r5$c4ct(�� �������ʠ�5"˦�����4���e<��%ھ!m��2��qG�m�eξ���xi�E���#^���������{�29?�����c�0m47i��O���G$& �a(q�v� �#��z	�� 3W,��,�����Γ�)M����ڛw�%kt���G�g���y>kUf��B����~Ra��\t�����	-e�wa �Y~�_ӥ������bsQ��x��ca_�xhx�4^�O9�@DgBXby@ �9kuo$��y�������V>���s�h-�c$�y�da�Dz��{���6Ǽ 
�)Ru��;��E��n�۴�ѐ;o�""2^WK�&gC=�˯c���~nvZ��h�d��E%s��g��ٝ�4+�҈�ތP���&��c��&b��߅2i~_\>�@^r��Q��9@x��qhx/��s׮5����VޜE��dC������rQQ��#<P���d0�=��y��<mv��V��0	!��9�T�5��~��e� �����2v.����o����m�VKJ� �>�>d��!|i�%\B����8:����4�L¤�`�qY�|�U�&��5
qXԾ7���']W�������m��7��&�%	��YE��y�̕�Og���]`՚��7��K.A0h6�- P5���Wu:�%�.|��l�e���ѭ���'��y(�N�t����I�|y�S�2R<v����w����: 
	��]K����O�Tf	'�����s�Qg�c$�T8暠RM�[����lM�O�鐔+�뎄}�B:�W$�U�ķ:Sh2�)\5��*�},���廓���Ax�H8��	零@H�%���2	�8�����]ɘs��/lD�6G&*���v�I��QuM	9D����W�-����Au �d���<���v��k[hN�]ބ
u�2a���\�H^�T���G���X�KK�6c&�n���\���'��,s��"�D�;l�^ ������K��u[��`S�\�1sϨ<z9�I���h6��z�Z�5�PP̰O��uPx|I�*�Ov��|��+�}/�8��q�o[5!D��b�<0í(.��[r�I8�4x/��Y��񟠐ɣ�Zd��t-]���˘ՔrQP�>�.�o���>m׷K��L����(y d�������u@T�����X���u�?��G��x��ǅ�k�#Y�/9�t��������a«�Ϝw.:`�H����D�`�=��g�j�'H��.�T_]Z���f��"���kps�LY!q�I����Τ�����#畹1��E����l%*FA�.�ǧW'y�殟�P�Z�Uu׹����<��ec�A���x��n�|O�z��X�8��]jՙ�k"몋�g��~L��w-��1?�=�,�;�,����y�g�_&���A%0J������d��\SЛ?��{MJ��M'
j����:Y��6g�UW  ��8_���	��ܜI�@U���D
$;���C�5b��bMv&sʴKl:c��8x/�CPw ��h${�|G?����"l�u����o������#�BN���A�S�E���e�-�!dgO�T�:����	Zl�9@$>�(�0��
D!���ql���Gp�$_�� ��(T4����Bb�E�C:k�H@��v[NVG`� #��Gd�(���o��c���"-�B���튾�z����g���;�s��5��h�Vʍv��d�<��2sD!�eFXÔ��הP�b�Կ�/�:U�L�*�T��#0�o�H���ݠ�iDJ�[�Jl+vO���5w-�T�$ ��e: 57���6?���5��h=Nt�I�7p�W;P���x��EA[�F����%'=$OkS�X�0��v�B���M\2mc��[���<������m1�U&�����H�+1��nt*���J����Q����j����z�mY�ԕ��x�Q���������fѲ�@u�&u�P&Y�°��{���H�6Y�e�Q�Y��!!�Q��z�x)�l4��)���͞�w^�`;�50si�im�<�$ga.��`uQUR�����~"��$��_�']��ݾ;,�N���6{i�r����5��
��%�5����lz���$�&^�^���e��0���tx�2��x���W&����!]����[<F�kI1�U�����.��*r��q��EMA�T�R�� �<7��-xQ�t���`"�Kv���U��)�N�(.`��~��Y��T��u׻��.�Ce���%#dvO���Gqf{H��f#;@|F�WT��	
%���Jv'z�3�x�"De���oR�>��{��b b�tfה����A+H�	;�JY�ΰO�]� ��LU�mHA�H�ؕ�ć>�9�=g��)vr�@��q^UW~��@R��U����\ƲCǠ����t��265)���/������g�3f�>�����Sx�!v��l��𽋞 (��j̏ġ7��o:8� �\�5 �O;+�����w���J@�p��OþON�x��h�Y8B�t���?��U�!oqi�5��Vu@%��J:��A�VP���g�3&�qT(�s���c�"�i^<�?����a␨�zu�vv)�w�m��r�2����Wv��@ Jb~P8L�ŷ�����	��̍T��J}��]Z�_�+{�6L����Sa�ܠC��ki��m�羨�8�(9uRj��j:m]���3-]�ӑv���ͺ��fXn��)�I�̹^�����^��V`?Hj��'��iе�g��WJ�0\o���$��*w�/_ڻ�	O3R�牟|��g���W(Z�P��<e��^�ն�u�
���<�JO�H�~�%���R�����x��_O]�a�**z���
l�q�PC���γ#��)q��B5 ^� ���v��6�^巵��a�'���J�
 Z�'�x��K�����rwG��[�4��7��}�I&���Sވj��-y�1��|7�t�JI����χF���z�����b�"�߯��zPF��<ψ�:��O�%E��	<^v�'B_%�<1�B�O^��	�����g�K�ڑt"H8�\��q?�����~=%:%�`��z����ϡ��E%�������v<~�`�T	���fm��Oc5�I���z��V|�ҧ�^���Aʾ>����}g�+��g�⋀҆���|�g�����g( +Es��k������np<i�l���}��<I�
�nu� �7GI��JX&��I;F��D���sF*b�Ƅ��䮏
�}�z'{A���6(���:/I��ovd�Z��Bsq�֘�/�%������*�@�-5ξ��ċ��|6���d�;A���dd�IWBRmO�1%���v�K�Ho4u��hT�yu���3��`��r���y`gӶ��L�����'*8���O�[T��ۺ�R�
��hܫg��SA�^st�3�4�|-+����X�qԽ�Ҍ}"`�Ϸ��]�E6�4�8{�΃�$��.������
�&Q��=�wz�c�[�����ʢ3��Ы'F�BJ��.n�"`c�Df���r2�Obi�8����0�yL֣�+3A�;=�z�tu��r��@�&��&{,Q��ΨM����w+(^�.��hh�,�DۚD$�P��bp��ty��l�r�t��dq<S�x{9zB�;K��^.*�f0�&���@��� ���ҋT��S��Ɣ�+댝�[�i�WO��,D�Y�>O��J�i��������w�<2�dq�L�{w!���En@H�b�����
]�o��j����J�PR�.�򴺬�]s7��#m�wЪ��]+��	����I�4#�sr��c��32�Q!:B���d��Ʒ�������ˍ	�H�C��jw�a�Po|n˥�nҭiنj���K�|����uuƄkR��!�!��l�:Ґn�.��Mf׶wxQ�.yz���y��Z��=1����U
=�z�#�~1'��\�wW����V��2\}�K5s=� )Xck|G�*L3��moWٕ�ix�?a��P5��	�/��oH��<�l�a�kL�츥+]��F(��j���?���]98X�?#�oD��Y�L�����DrQ�2H�y��,���/����la@6��B�E�����2[��\���>ꎹ��7}x�O�2��A�ʍG�aoў����սL��G�[���'����j���B���s���cV*�|'9u�T���0��e��s��ͥ��x36��Ǣ��W�
�.ɹL$�������y���(�<�>IUp�n�2.W?<,J��~2���w@;���y�v�,M��buC����Y`��o�{�#����-[�o�%(��,m��譜���L<������^=	F��܅����������mav9��bj{�=		���6Z(ՋEE����24Cވ�$9K|�.4n�zua�yl϶��9j������y���Ӯ�ԡ�gR[���T�s�������h [��#/nK���s�uHK��0t��wd�%b�Ou]/,��Ln�2Qޢ%�玗.��#���msmh���v��:Q��-J�S]ؤhl����q~F ��BU"ř���}�ku��@V�kN���u����ޞmq9C��r��uG����t*�S�Q���l��L6!��;����� ����C�V����B�����~�#Ui�����oM`[�=#�̱ ���1�E�qi��t@�#%���QaP����Q!�GG% ����0C	�~���ܿ�>��od��ʻ޵v	�"�zV��FewR��h�|����]������l�v��}h��S��N��N�}! ��+Ӡ�&�y��ǭ�t�~Oi�a��3Bҝ[\�K	���a߿���������"���Vg�j9��/I{�+�s����/��O�5L7p�Y����g�9��m�������ӝ��ޜ�#�H	i�$�46W�������wt�\���/I'QFF2
Z�M�p�֐������g����p']ϓ�^]y=�lc|7�ǥ ��ش����~�Ѝ#���,���F���*ճl��1����՟hY x��};���q�N~X�<\��T<�t�a�)9*���f$��{�CR>���sq?�ɳSV��\1��-�ҙwa��V͹aFh}���������P��yqR>H��6pW�O�|׍�0(�> ]ڄ�"�����A�u�n?�ߩְ�ʼ#�t#Ь�)Tf�	�x���+�g#�sV���x0��Cr`�"�&��'V6��cg
�.3��o�A4��� A6��.��'o1�Lذ�⊭~۱ޑe����;��
�5�����'��VHhQ�Ph�>Zl��q0� I(�la�B�G�o
�*;xtwoL��1@�1��^t�l ����*��
`Q�� ;Z��?G��EF�\��m]�+9�2��o1n>��H'b��/g٘+ndn1�9:\]�[���񤤰}�VxKNI�K��w� (��uC��-�Z��@j:x�񈮼�1Yk{jgs�mip ��/%�w9�[#ۮ�f����a�& ��駚�����2?�Z'_��|8�)Y� �����P,���t@JhrW��A�7!b�
���o3]�������ʺ7>����^|I�[�v�����n�6~Ǒr�7=݇�2�?@�����#���m�{��
���j�I���p|_@%]�:T6� ������K�Ev�A��+�y����U���y;�hZ9� �0d���~3U>G����"�
�5Hm�%�F��������G�����ĔU
��4j�mo֐��2�`?'����	�i�\���3�bUS=�K_�}�
m	o}��@����O�h��`�ʦ\�����L
�&�����#������������"�[�_@��Ji�&'�}���)�x����?�01W�r�4��O6HS�6�c���|�^�o�9�!�X�T�@�!�!��� ��M�V[�j�'h20E�N�*:c.�᱉eJb�~��yހ?1�)������u�2��.���34c�aÃ����n��9��g�Zmo��� �{+lO�ģ����&�ʁ���i/��'��q�*AYR_֟;�c(�D's��C�x$�M�4(��h���6Yk[8��
U���^�F��`���a������l�BW�/ut��M����̛<�?q�*���Je��ﴞ��!A����]�q(%	� �%%�R�I�ہ�&�4�������}Ru���9rG��|�KIA	G�zk^�A���$f(k	A��gx�W�� �����ZSۚWLr=@b������ �퍓ɂ�jI�?)��>��_�w�1ĬF�h��Auhn��a����\(%�	hvK��v$��@3�+u=��.(i.�;�b�>���UQK�:R^d���o�ȁ,�f�i7p0��c�x��`K+�kO�>v���j�
�Uɸ�t}���_��R�D}GA-
FWo
�
�1^ �ڟ>"lQ���������4jr�UT#x8��8J�-Zp�xv@m�_W@���)����-�̜A�æ�ӱ0jw��9�bW��`��Eࣀ<*�W��-ț���w ߗ���=}J I����;��y�e�}��f���ap� p
�6�!��lO�⏧���C��H��)���X�Q`_m��_��+���6�w/M]0J��`EΙ�Ԛ�`�l��;��g�A�\�f�9/�����Zh���)�W�7���رƈ�7vp�M����,K� �����] "R��?�������^rV�T�F���"�{A/�:(����\���	��Ȧ�N#{�N~�X|E�yʦBi��E1���f7jy�����O3���G��y�YV?�66�O2sO
�����-�H�c��!u��B��V�=�5+�6�ݘY�W�����c�Xv�&*�A�v��U.r���폚]�7Lpo�i����k�mڳͳ�)#ߢszv�j�� ;��HҀkYpc�|J�w�G]$[?b*�o���"_:���Xۡ�9�1�7��-o�����	��k��<E8�E�#�O�}��������+�Шm�r	��Ja�e�I�ԶYmYZ�4��R��)��B���^ZB��t��4��ݔ^�)�$`O9���#j�㖛��N�E;3~Vhw�+ħj�y����r�ޭ.��j��2�������O��C؂�IU�jo��fVH�l����OqLo���tр�ᨣ'�d��#
ծb�P��������++'�7q?
{E1�h}]� �#>�G�Q�=���+{BTM�zK%���jӋ�qڍ7���	�>|�
���4@d���
p=�l}�j_�Hm�˛;�R�z���RÞ$WS�E�@	�G�b;�j�s�o���5A�,��V���4��˔#�?t��l�@)�Pk�:t�Ӑ9�-�[(�'Wa��q������{Q+��.�����Z�Ŧ������(-i���[<��IQ@��iT7�h���Zv��3?
L����y�8�#G�L�쉩�
���2��A��y��#�̋s�b�`��^������	��r����ڨn91��]�i�8W���l,�>An�,��8t�\�]�Q��'!D�C��a��Q�.bl��kLO	�)-�S^P�WnEXD���t�mw�H������r�i(a��:K}���R�)*�T
;�J���%Wc��HDy9�.���H#�l�N~���ԍ�W����-��[��R��9VD�����>5f��`W�G%�|{Brr�\�S�"%f)bm:#���(旿y�t��wMsB�}H�ǖ��+lQ'���ز���7�\�	=�V�	����vͪ���Q��l��c����J7>$n����0B���nbF�Tj�a;�iޛ�cիGKo�b�־ƺS��������H㦨a����n��u���_m�k�<�j.�1xi�d��O�o}T�b~�B}e�L���DG����P��]zQ7mb�t���6o��2.���?�4S[�<cɅ\�G�����o��_�a��Dr_QvC+]Gu�3�}K #�\��Ʌxëo��q���Z6h�gr0��ϽԨ��3�{7�\��lsh��0�4�y�;�VN���@������P�7V���N��kf�fpc��p�rխ�K�����D��oR�,f����d��;'}��гue��Q�a`�b�������x�`���^U-1~�ϰ�Ϳ�]W��Q�j��kO/.�};4(8�j�0�]��(��y��'[]���y��|�m���I2h.���	?�B��/,0�t˸�$3���O�~�)�63�W�S�i�a�'�&Ҋ���we�MJg���ʩKT�<W1Z����W΃j''�gf�M~���rz8̞hg�c/��.V�����y`�c�7Cmߢ�|Æ����V����P.Q5�K�:������I�:�
3��q��۠g
���J��Tcr�z��*��Q����baK�,<l=����鄟��a<�q����k�i���ư�W��T	����@�$��4$��. ��N%�s��$w�#��4�3��7r����đ�d��p�
�gF.�%�p�D8��b��%uz�b��d�G䄚��`-~�=%�ɪ��~�u��Ah<SF���On�B)2��%�7��g�Î�@0�Vr��o$94dbw=3	W�ݤ@�%���ri�)�c��:�XI�w�����=��q����J�ѺW!X���IYY�ۂ�\�Ny9�t��)8-#>�G��:Vnm6/�{�J̛�|�D'�CUjR��;�����aL�a�q�ϫ�ʲ늱"�BIFi)����*��F�Gӌy���S���,o
B�w������%mKS3yRBڟ�v�^T�v��T-&E�V<.cf̭�u�bw���T��x+���"�d�*%�i�ﾓ)� �<b��x�ՙ0-%����tfTcFv�X���Џ$tx�Ҡ��&�ha������Č3	� rc�ٍXL�B�*�Ж^?�G>~^��������(������P�O
r$�M�?oa� Z�)i���������$OPޒ��(#�;!I�P�9M��Y�/���B���'��N�^zq�S!=_J��߲o]5d5�h���U�3:Vݵ��<c�Tۛ�,��S��0IZD������xl� �j�^G��{�PW[��\r�Qn�%��O~V��*4A�d����2J�#f$xv�,E-դb�#�5|rD�'ޠx��n��>�b)���NT�p1Z��B\���')׎D/�k85v/�?l�Zr�����&�,��KJ	��֭D+�ː;���$�骐s6X�l�2:�s�N�Va�!�W\LD �U�{��7 +��aY�P!��gH�(��3��B�}���XIfaw�T�3�+73���cBe��UЅ��͵���f gj�Pb�_ס�%
��v�h�1�O�37���r��YU�7��O��	�MQ;"Ͼ�N������_��*��pT��{�n���9t�8)�4��%��n����~+-�h���`���g^hD$�(+�^g�j��7��8�J	�y�F:4����ʠ*�uKq�j���Pp�k!�!��x&+"zג���K>d�U�h��~��#6��<;��`F4��Y+��G��%�.�9��M�PK�s��ߍ��d�'���֡.cH^yk}�����T�9�IVr�{��y$��k/eH �]��.��
��pEe�	�k���q2��sB�꼚p�H�ctONg��DF�>�P�]�q�QG��z���BE�!�	��]�İ�>%K����K��H�J�x�憚58��x��W���H�R�@��	ڦ���|����#�͂�=��?���5�$a��fV��@�	��մ'���kk���'��z���dL
y9�p��N2`�b��0X7Lu �ȱBzӵT=p����@ّ�P�&ߩ� ����ޞ�k��M7��8��F��BM4���6�X��y�Tz�4~ܾ:��F�>�	a:c�۝�a�o�>,@��'1�h-^}�h����z��&�$p���=�Dޛ*���%�]Q�b�C7e�0*6ϯgE�����P	���V(����0�=��M3�DP����k�T`�/)�Z�J�(e�������Fr������W��Z��p�q��0�y��ʯUv��se״���V��ई���Խ�!�g��e4s-�\�����4z�K�qU��s��aĭ��ˢK1>TǛt�i�'��kLҰ{Q����iLr/��9�o�����Z�A�|U��~��|8=�[O/�C�J�r=}�����qMJ����z-V u5@��U��FF5��F�Y�F�bL@�LX=��kl�ə�s�	�о��|�`�����t����pB~�%�J�Bkw��选n�U���d݉2����b���ѐ'ʸ6C!v$���k���SSח������T�N�>m�:�f��T���K�:���+p�Ľ�ļg|�R)��������V�ժ���՜�ݡ��?��[�CTz�a��Q�KYҳn/�2LY����w��R��B��
?�#K����֞ľN
��$3�:}6�}��;����?<-h����[ jQ��v�OR�k��G�����$/���|�ӈ���ѹ���&M���|��{7�T,���Ҕ�'��=~��ݹ��*�S}L6��Bӵr�/��$'9r�.SEH7��G��ń��/%h��	���xч؉�y,�&��0�Vr/s��Wd˻�n�pi�S����\�"K/*��p��1�� E��z������C�B~;�B�Իs�N�H��T���>i�]?�c�Z�a69]����Q6�M��:f`�Ϝ?���A{G����E���|�����W6��MZ7p�"�f/�i�`n!�'w�h�>�g�I�R�I��A]�d9g���欉��Q.��|���4�:��`�R�����Z�T��<�(�/���S���4����K�JHF����^N1Q��5�.ũ�*�����[+�ֳ-*�!+�6&2���ˋ�-j��}ЬXFc��ఁ�β�Ɂ��_�����a/�H�N�c2B�Q��	'S���}�����I�=m�V�w������ڠ��_��6T�����q��S��3p`���^`�L}�+Hd>��Z��B��Z��AD>��Od����ηxm�M�\��$lO�m�K����F�F��h��7J�u�90�l�*C�9��+�J�����=0tN�)6���6��Cp���#n�ژ��{TB�/*�"��x��y���e��.�YWr�Xⳙs��aqȺU�dE�T*��!/N����lav���� �[�����g����Ճz�m#?� Q<+������L�JpwY�ꠉ���w�(�r�k]7*�Vꞛȹ{��iቆFl���W�$͹xx���������:<�VJ�=�}���ӟۤ���{�R��a@:��OcCG��y����	�3d4�S��\O�/Q=����a�y�|҄�|�0/Flm�k=�Zz$���0|���d��f~
3y��E�C�b㓅ir���n�uĘ�R6����o#�����ǧ���dv�EXB�qH�{u����CGӑ쵈#��~��NL�'���w��9꽐u�܊^#q�S��J�,(�b�T��������&�L]���W�N�t�N���-8��+7	׿`��+y�w��>#X�&�?7�X��(�m�GY!C��z0A���+x�~������8�'[:BV��u�<�t����v��F��-�'����-������y�4�R�z����8���-!Z��I߾�?'3RFV�CU�ӊejQ9|	���
�C�7q�r��a�Wߣ}�k١<�ƃpMu���%ևu��͏~���y�ԫ�����`�����U����
��Q��I5��@;��"���d?�m�z 1��&
Y��w��� t���d�e�IɎ�&��"��'��m���w�2+܆�.#"���@��5��#�!�gf�aiʻ��0��ޮ�߉�����]8��)��׆LF;�̩Ӭ,Z#�����{��g]�����{��8J��-�����δ�(^y�A�8�?�j�^����	��>5�)ړ- �lp��>�wv[�����x�8%B�s�O��6R#�s�;�͘{�ZS�<�HqpБ���to{s���`�Od�t���(��P� ]Uq]���+�^�̖����_�|S�x+�)>Qx�K#2^,:��=�� |y�0��K�ׄ��'��kC�����Ҋt���x�ʘ��͈G����wa^t���[�1��N�d���!�CR���]�����Cq8�;֟$��X��d�QE���(������
���lzn�.��Q)�~�5_;��R�E�57��ӑ+Vl(�C:��������Q���W�-�XTu��SF�$f|D�ch�/[RyJ�.]�����z�G7��u�-A}T�"�H|����+����ۧ��:���ď��t��#M�
��5Ecs#vrP6=a�6�E.Q�!X��c��1���pHM-	�ĶsD�M�:uN���L��������,w�K���k��[�z=b��~#�;r��e���t�δ�5|ڣlT+��<����h0��T�.�-rԳ@yՈ�F�6���z��	Õ䄿�o��]:�L�q^��Hk�s�k/�����'�Wk��q���KGk{���6��=܉�/7����Z�ӝ�PK   `��X��НR5 �� /   images/52cc771c-8bcb-4758-820d-da79c3626c72.png�uT���>:��GApD�tH�CiP�D��;���i$����;��A�;�c��3|������οg���zY����{?���u_�u=C�e�����@��r�з AĨ���/�eo��[ί���|y�c \�u��v��~�~n4[�S�H�"��fo�7r2��pN+;��������E�(�$}��=ic�#$�؇��o?�W,i��O���I2�j��(2���qS�a2-�"ؘ�*���AS�I�ԋ�TV����/�����J�ߦ����� .�����������N����ÿ�/�׋�9��>�mP�t� b�������׏�4���+�$n��x��p�?w�ƃ��T����T����?S�oSY����&KV�M���"E�����b�����	������KJ�y0�p�_��3E�~�@Ҿ���@�g8,��?����������ۖ/SZ���+]be-�sQ��d"��AǑ�����f���\X�Mq����U� f ����h��h<�G���U�,l違��۫2\f(.'FK�npo�ד��!����z�@mU{,)����&�/IK��#`�z���Z��A�?.���c�KN�*��}������������_O���.n�sOX^Zm*s�uzc�N.��:)�5J���<Z�`�\���wR08�,�9��J=ux
�}�T��	�j��s�:$�!��u �Jl��)����u/����_ f�m�3�!�K����@����އf��S�ͪ��/�T��R�]�_yb��[��u�(Ij�CJ˭���]?]}�4��G�zE(���]Ә���4Q�,� �ި���'5T�iy����L2���jbeg�VC.�2z*C�����8�\��$q����o��T���a9����O&���
�jVk��4�����z��q�P�㽵�8�u�Uo?�*-�M5Lz=n�s��҄ bW:k~�D��Z\}L��nxm���Y>����g�h�:i��5��w/t��s�*����3V��ʖ(0&�����U�_�W�5T��TSv���w��ް:�xyS�ˡ��Gc[��6�&8:�`����ӧ�ri�����u/�Mz�+o~zj�vTM��9<����x�PG�!�A^!T�R�>&7��p�i0.A����i�����ш-J� !�9v\����� A���J�j���c�T���ݭ_-* qNXhI�r���R4�z �.&09��AA��m$o���ȅ(��d@Э9#O+�y�`	�%r��.���l���ӖǪ�|����R��lߑrա�T��ʁ��,�k(���$�٭���UOˑ���W.�ɻ��@���|���w�U)Rpt��}E9�d?aqi#�G�唻��^[��(�L�^J�/!A�G\!�:��v�FaR�ա���A�������7��1�؄�q���z���x�3P6�?A���]�|5WD����k4�0))�$%�- ��t�cI{��R|��h��/(��t{V���?1V���0�܌!�RȓyeK��yV�n�O��*��5M"<u?��2����i���b���X���#y܌+���b�5�1�&9��N�>���F6~=��,��"���sn9��$b�&�f�&��H����45�4Z#��2������/�w�{�/P�8<�Lz��4z��)�\.��={�˷ O�ӊY�M.aČ�x��n7᠍����)�^'��՗I�5o�x�5Gm�GYr���:�_�n���Mi-�q���V3i/`3��Vlڗj9=K���S�;h{p���L��k��&���D����;s�?F��~�+L�t�X���<�6b-�l��Q'���s�$���c�k�0L�x����x;�����yı����2d���2J�/�=/�=��0��773x���O���I�e �{�ol�L��9-��	�K�+���1��Q*)}��F�蚍M�5Ml�|����=k��������%�^>6^IU+�F7X��?�cޤ>4�Eb��(xT�@�tf����&VC��Ӝm|��sn���/��j�p���B.<�����ȥ��	��C��0d���]�{Ι2��ȳ#H�%�:B�E|��|����{>�ф�(�_na#������^��oܹ%�*.��oH�U�O̙B
l#H"�wb4)�4��b���a�����0�\��:��Ւ���W]�����3�L��P!Lr-�|�}gL��+�����h��V��PM�@3���=�tcCV�V�{�F��A_�Q@F�p���a-���Q��n�z�O���7ۂ:>R��K�8�O2S�lD���׺�ǻ��Kf1���k��Ή��݋��2�#��^����`�S�E16�����	���T	�h�#|� I^��:Q�zGG�IWV[�'а>�0d�fK<������3��,�݉3)raĹ~�>Nv޼��ո/7.3�ں�N��0�{�C�D>��E���or�DV3��1�'(ԾV�!�N5D���}rjƵN*r$��w|�3�>��P'�=p\Xb ���TR�<���~I�|�<�S5�&���oK |��̬��"�jk\�d7O"�Q�4����G�w+��7M� �$&�?��x-�FǺ���F=h	��lRN�����r�3�y_��Pƿ�������ܱzG�:��)Y�Ǔ[g��^#m:0t��Q��Eiح%E��T�������M�D� ��E��#A�U6��U�h�vP"%|�ߵUԎ�P�r��4P�O�������^*G��⎩9-�-�P䳛�~Uu����1t�A��y{���|�C+�[��(����7衳�Nr������"�wۏD��\��p���G�ʂT�,#\�[Q�$��h�
�����%P��f�_�P�J�������T>Ր86ϟ*� $�aR�Gr��mR�n��� �\���i��p��Lj�9US���i�4:�,?��6�����a������MWq�x`1�fJ�|�6����}Hd���s\_Gq�-6�	����L��3���4��ب1���(K�)�&_X��^��;Y��wI��6��ji��%Ƭa�∿�G0���"��R����g�ｅJ�E�	�y]��(-�I���h�`u�{���~x���F�������2�D`�D��^WߢJ}�Q�H���M����*�nN��[Q�0�c/���}��ߩ�p�-t-��jj�TԎ��2����n:# �?�%�6�_�|�h�~>�F���m�'&V�-3��N�Vư;a�n%\!"�H��7��Q);������S��S�����|��;>���Kt�	`3쎎N�Gx!@�Ky�&�m�d����������*�*���B��vh�h����o4%(�,/zRPжY'��=k����9*�3g���"��׻"��'�Q��0�? Kb�b�
8ZX�ƌ��(���G�2Ι<#�W��b*>g(p��z�c���A��O".�!F�)�@���5JJz^!Z� P��]\�;�!�f��NW ^�`=�X�Jg���K�U�ll���#l���\�x�URh�}�+ٸ�����֦���?���0�o�4[�qT����cM�!��7����|�,:��$���*�����(bt��R�w���+у�G����tn�.朏�mxۏ7k9���`t�Ph
@�go���Z���*��� \��N�,G���������g���]�0��+�������	okϳ�0<�op��Re[��d��~r�B�j��Y]ip)�r��-R�!�X��K�	:����m��Bj�,Y��r��=��������Oe�S���-�����Xs��U�w�^V��oRe����V)��)�O�vfa����¶��~�ʖ���2F4kEa2�ULD�)H�Gs�.#m��	�'|oQ�@O{�A����*�V�t=�+9��Q[�LM��n� ��K�n�۲6����. �<����y�w��l-j���Q0�^g{3Z|��A��E�*�3�< U�� ��R\�?����[�� �"�g>k����&�M z[��vp�䂤H:�nw�lOq[���\�g�������G����H�.
Y�C|��	�ު}�,�¶j��?jk��z��
����O)>�>�� <n;$H�,|��j5��z����k����0 ���l����CA��U�I�n�pw�Е���6�E\���s��[W����<?��=�7?���8V��u��zW���5�r���c&�q@���}����^�@z��ځ��)�m��V�S4|��ʲ¿�]�ud�E3��k;�R�;���j@�p��Wa�G@�\�1��aT4��hK'�zX_��-�a�#p�#�T���(�qWa�²i��uo^W\�Y�>�[��0����#��kp���~۷8��� p�H� ��}�SN��6_d(�����]���͐�Ҝ�}��y��
�]���5V�oܒ��Gn�_ɍa�!@��/F࿐Q�TQ5�H&�]�n�D�H Nj1bv�t�(�#�}���ΘIp���v<N8L2�\���Wd�-<?����yk&;����W�_S�;0}d�&�0���+|�N���޲���Gղ�
�ݣu�v�㵜���:��!@`�Ϡ�,x܌O���Eϖ��aKD)C PZt`+�w�2��y!m�g�g��C�ne��)?�A��H�>z-?������+����K�n�e���&��ȍ�-u�.a��kd�P8h��JC��;��J�n��l%ƶ%S���r�Z·�7���>����
����J�����gQpƘ��nK���i�^�;ޖ��̭&5B�Ϻ�7Aa0d��J�%a7����}�@��03Qw��ׇ���m��]��,`�8�7��/�Vns�	*.[�W�K������-ӏ���[�&5́*)�6Iq��k1G?�����Q?*5��'M��-�_�>�c�h	C��M��Q=�5?�*���1��I��}S^>�6�/�*�3��C��3����i�qFO8*��>_�p8��o0�����ƻ��R�/x�N+ɕ��ǚk�va���#�s$���6�?���x�p{��}��� 2���}2W��]z��q,`���x�����L͖���x`�L@�ğt
�"ị;H������kP:��C��b�x�8�h�lf��L��{��ǚ��=�?���O)1���bk��%��� ��> ��VZ��nO�h��ZT�2���s�]�\l��y��a��^R���7K�����F�;:��,���\�,��gyl ������ �&��#�E�{b�/q5�@I�e�"-���!iriJQao�T����[�Q���G���V�.R�G�r�����X+���
�(F����[�w!V�Ph$����e�+U��	�{�`+��r&	Y�P�/N�s
ν�����\��D5g��AM�"�$�����f�g5_��e��Cr��Y��&�Q�L��+y_���V�+a��'��BN����թ�<���_=#���2BWe!��.��r�k	d��߈2��frQ1��DB�O��+���3=��
��;�U�ȟ�k��f�s��IdF�U(��ڒ,��`�	��s��T;�
&d9B�"+���Y�O��9դ�-�:���y%���c�)��D�/!��z�^0��2��1Ƒ��<L�|��f��&�z��NF��Rzc�c��%����
��xջ����H`�6�x��CJ��Y>�aN�V �d��ҋ���2L��-2ڣ��Yk�o[r^G&��.������Ọ�����;�$�͋]�(J9*%�'��qҼl����hi����F ���Ҟ��D�k���V-󀓖��)`璈�Jqm돡��e��t����`w]�Ƚ����$K&ݒ�C�2: ď�[K��CDZ?��U�6�w4���m����֚�-���|D*�������G�0H`�|II'0�l~���2�+�2!�8A�14+�aY��<�;k@�R��L����_ :o_IB�������+|����~!)�,ٌ����a��y�����W�>�� �(���;��`g.�?'�3�GZ�k�O��9�P,Jw���v�fSO�cs9�O;e�V����?� �q��j<�a����U���Ռ�c�_vޖɳ9V��h�!P�dsE�"=r�z���l�a�ҳ؉BJj����R��f/��RtU�����zV��6�
K`&���>Z���sC8�H��ƒ� ���%F0�3��I?��{2�IC3��$>�t�������ߎB%�
�s��V���¨�U���n)	�Y�z����6/h�
����YC[�����������u6���Nb��Ĺ}��fPN����Ģ����K�֮��u�����Y2}ip�A��S�.cv5���a��������d�"~yo��^������N����Vr��D�F'���������t�5�c�%��rz��[��)�㚓Q�:�臼��I)��盄XO_H���۪���$�o�v��=�>����D3V�e���@�*{ai;��� @��H��f�zA����)����)��-�nQ��hH��tDKbDF.�>2Q�C��rU$�q��G����u�!M�_?Tt\Q�zFԞV���|���w9�n���;�A�J�nN{�0�"(@ b���K�9���o���������g���

"�ZI=Q�ɔ+y�#+@�D���gCJf�+��O^6�Zg��}w%�o*������(
��͎_X�_͙4���֢%��è����V�?93E��ӳj��Y�+o������w�Κ�K�"�Z�k!		%a�rk�z<ص��0�,���l��)�!Ҋ���+�8 ���� oO��m�!�#�9r��E���%�Er<�����Kw]�]����!['���b̏p�"�$W,��$����Y��=A������gg֟�'|��B+��%�({��׫%���`���犀���HdyN�]�xTJ\�J�8�Sav��v�@�K EM'���Z ������*���BƁ�ȷ����K�)�.�zVjj�o��KX�
dM���r=j�	����oڹŵ� 1p1d�t����v�����K�!�C���6�e����,3ӭ�;�o���6�����0!R����x�pX����KZ~-:��+���N��*��j�w��E�>q�,%�jw�T�(����9��J���6�1;u��٫:��:��@a ��֎0�&#Z�#�ֹ-�%�k{��ә���t����p��v4��g���_�e�+ ]�xXc�-t��rs_�i@�;��h�:_k*�۠[Z�uԱ��gl��d����R������k7��2�ohTf-�xD���ki�����l]���PY�`Uз�3����Z��~�ZG����V����ٗ���V5�ƶP#[O�q��o S�KP�f��L��A �~�k.:���y"]���2

X zuD�8��g��R��$�JZ�BfF�T�;����l-��`m�΂�9��&��F��	O}����|���Жm���^�F���C��B,��BY��u��s|wGL.��(E�m�
��XE���㩓�ψnR�m����)�:;޾jn�r�2@�lcG��߳�G�:�F�J-�:6x�/�p����m|��pXf��x�hb�đ�q##�uY�h�H�ӋګAbe3��h����1xw��bӞ����n ��Ӟ�؝\6�K|w���8�EEqq+���
l/C��lx �nߖ����ɨ9o��R����+��6�Q�-�H�o�
VMQ�&�:���k�p/JK���@m؊r=y�~�a��Ү�)1��QKC���h��?�F ���ϔ��	�LXA�8
 �K�)� J(��֠�/���H�\-�c�}.f�,�
�8���#]ӰV¾�[�E*2���?��4�j�)��&H�S$�6@=�X��0��-Z���}��rgE������d�����"��h����y��xQ%t��`�Q�v�(���m���+�Q __�N,}��ta=P6��$"���pC���}���-����F_&�(`0�g��.fE�����J|��Ք]�.�N;YW��O{��1��mL�_�Zwڔ ��׽.k�������/�����+q�mPC(+���^rHK���} �%)���Y�у~Z��l2tm|/!�B4�zA^9Y�LlP��<[���8�,7N�)+�a&�b��t���\�8�L���﬇����b7[g��N.�<��m��ϧ������υ�N-u��6��{���X3Z徤�����n���Bj����qt��E�l�]Q�.{.OjW����bC��Fp����VC���&��XX�ǩ�q�����%��~b��:��p@W�d�6�I�cR��Cb��W���Z	J��BHi�~l�v��Ka�}�JA��@Q�?p&`���͓��eR�>�D��1�0�V����PoH���F�r�@�B�l�x��`�^����"��٦2X������7c��$'�jA��g�i�#L٬ˉ΀3�MQ��!�՜@
�׏�$I}}G�H6e0����B	��s0x7���c��v?ĸw��D���{5K��hO��u,�nL���l����| ǧZ�Y���j�����ȸoݖ�hc�y-�e%��i��ޫ�˽픐��}�e&m��Y1!����4Tx��i�2�12Jut<���z�l5�6���,䆠���h�����;�T�*��xU\lw^)^_U_�P˲����/tc���އ}]�E�mm	�_(~��3�{�g�\��B��Ӓ;��j���Լ<&{	�"�0 �!�A?�7�x/>s�&Ch
��Rq���ZFA�H�7{'��X�E��h�Z�
��H�zZ0v�װ!7A����S�/����`��U^$��la�$Q�1y���g�Щ�M�1�>�������)�)-��$i��hBբ}%�n�~X.]���o����U!g�w5�$1\:ɳ����d��y�Ss
	�{���秬���w�L"a��˩����N��ƭq�����iO��w?C��Ro��9w����G�Bd�}`���O��ｍ&�� �f~��Q���O�=���K|����W�ܢ���+�+���n�/bCw*�:��_�FP�ǲ�����H:#�1����j�st����Nd�_�$�$�a�,@�ݽ�њ){�>OҽR5��mw��Q����Z2��2�B.����S�X�#y�r?>f��wj����|>��a���&P��@c$�Ux��`�|��{pM�`�i�eeA�Ƌ���*�	�15h9�0�&���w,��$�Qo4'�yYV/%`���N�d�2�u�f`�Ŷ��ö����I�s4yl'�CD�T�Q���1T�l�;�h ��?���E5IQ�6f�c"�n�w�i)�<�QKEm�xrE���2a�ecP�2��jX�ƽ1��=�9k�THJ��l�*�-�bX�Ҳ6 ��gA�����Y�m%�n�����0|��e��� �	2)�$jh��+��ɠ�l������Ѐ6���zV��
:��{&�;D7�AM)�E�:~A��>�z4�-�-ǸY�VTn<��ZrA�.��#r#ƴ!n� ~V�Л#_�_ޘ�r�!w�q���5|�\[�^�^؈�L�u�=��k�'�`��pe��
�[�X&����+��O{�я�}t��!1�=�}c�"�v�bln���3��j�a����`�˖/�?lt�'��'�a�N���a����~��:�)!�b�o{ϸ��`[5��<XQ}J��׈7��<�H�R,b�|x�R���p7ϴ���\z3�b�kʄh�3}�C��8�>J>4�#��������c�mO�UK�S��g��}�	�@���mȱ�QU��"w'�f9!�:AS�2:�qΡ�l+����Ǝ�f S��N'ZoЋ��·f��v�5^�Σ���L��R[�њTi��[R�v�b~�EW�K�g�����Y���ղȾE�׀��'�r�Vy���������"K���`I^w���'񄋦�5����S���B��n�T��B�m��.��虚��m=��:�E3�}���{���{m)u?�7A�.�p��o�n>i��OJ��M�L)�l��#;�2+(=-#{R�>҈t)�,��Co�A�֡SV{�"J��FP���*�jK)��hz���sH���2)��T�CX���W���k�ݻ����VR�;��N��m�����Z/s�A����*�#��w�İl�^pq�w>�!b���3�������6b3,q�2[}T�Z����nP4�?\A�����7{�h�Z��B�x�%���w*�K{�ߺL�t�Y h��d��u�7�q���fV��@�yG�\^o���=��3<��'�MQ�d&�C��໒˼sEy��d�j]('��_����Hc8b��ԥrzхפ^�ѣ��A��֊��c_��&eDR���A�N�.���ͥ �ZZS>	�)w��~��o�͐��c��ӵA�G��>���{���m|�c�`h����@�A�����!־��e�y!αH[��)q�����I7���D��;>	Mp������o#��LZ�j"&]v+��ѳ%��
S�&�
�`+h�(����/[����7��g�/d������uPt��V��Wb����W��;��jA?�>���a���&S�7�vaͣo33!}�B�˾���L>���2ϰC�'|@ �+N�(�Fy�V'�{�ٚ�I8�>Dk�.���JM�E'�����9�#~�ƶĦA�J�Ge-Й�.��ޯ���=����}�����]�E�N��`�X���U1��¤��Ԛ����F/nSe���i<����x���u�yDx͞��ή�wOJ���+
�c��ӓR����#h��\��uT�l�4�q�|l���~-���eh%%~�[փ��8Q��TUx���:�<�-��:c]v�����b&U�z������4�L�s�t�ߧ{�;9��x\�`H�̖�n��� 9�mYo�h-�=�~MfV���K�
���I�5��9ƦC�ώwhƿ��[-����h��b��o}���cؾ�+ezb:u����ϟi`��$�.�Eh�����PX㚌��q���x�����ՠ�9��PT��D5Dwլ���heJ1��$�%UR�ZK~�`����IG���U�[	��I��f	>V�?����Ͷ;l6�E��KpI�Y�o���5�p����ﲹ�30�1ש9s���*��n�׏��$U��gY����c��xc���5��e[�**i���[��k����-L��Bu�\T�:��Z�Q�xi9��Xd^@�s���N�,��5�I ��7O�̻_k1�н'4A	5q���q�8�vc]~�LT�@�p{��������I������/���L�kA��i9����l�V��t� $:�-��C���Υ��p}7A3��_=-=T<N�!���K�����]��y6�
׶u]�������F�)��z2���YZ�@�~f�L������P��B10�H��`w�K���v����	�)W͙�,R��>����Q�Eܩß�Od�o����E�����!=��X6�7P���&+W懗��%���n9z��V@~���:j�C��\j��Aְ��Xx�{���)�� ]��ȱX҄]$���Ɲ�(�(��5������M.�d�_C��� ���[e#�TDW�~�C�{��y&�(ө��Mr��#/��8u�g&9�8�?Xv����FIun����~�|�ψ~E���S��7��-��6K������ޅnwv4�I���ª{i%ֳL=��)%j���^z����Y�t�͞A U3���k�p�?p/�����٠7��j�)|[	>]�DD�tx�;��/L� u��W��oݞ����(*(xKBx�-PF�}d�uC����@^s��1]��EH�5��_���mQ��,���z��X�Y��M����?��_��Jߒm�C}{�=O�e򾥽@qL�-6�6.QO0-[�,[i�7���Il�TM9=��3:`�.I��6,���nҞf�F_p>�̆��Ӈ��[Uf�=�cEڞ]��m�/q�=�R�Q�]��`[���׆�*���.~xK�2�ga�x�U0F�a��r��h����a�<:[l�Q��c&?��)�>��0�cj�h|Q�FM8���y��OPFu�O�4l.�Y
mU�ۏm�N�)�I��I��>�|ϫ �wR�D���P��<]G�	O9�OΚVEi̞-���9?��&��X�R��b�D���g�ު\�/aX�7�X)�.��'�?�Zk-�\+(I�|����\f&��w`$�~%/���R���%����c����(�ĳ�r�1s�	�΍~�!Vӌ�q��S��9Ǆ���:0yq��M���
�`"j;m�O���_.�<�pX�ѳW	�:�h�����-rd��N9%�'hD��b����:��n}A��(e"�N>>z&k���ϊ�"&o9�9�\����%k� �S��^T&��P�����X=U[��Ng�@�OFs�=�Kt3�i�B�e2NH��[*�׏w�sD?��Z:z_�5�-�n��%�{jZaC���Vybt"]|�����*ذ�"���9���q~�^!A��NcX�żW���!�e��4v�Y�/�K�H�א���¸w�����m�l7����į�/z�*!��J�8N�35��ŧ;�\�S#n�V@/��$���!N"|^T&G�|R�u����q�$����A�V��Dǈ��V�c`7n�[��P�΀�xe2�;}��(�ֿ�����h��W� �=_��ӄ��xF��"_ګ^�%Bx��M�0=a���Q�lNE&����H�᭦ᕑ��_��Dn��~�����[s9��K�l�����Z^��q�D%f���%�e�[��>�I�_��\yǿ/���=1��cb�Xm�,�_5����3uP���7�83�uTK*}d�W��/p|�6��/y�˳'�Ю����gO�m�q�����~VA�Z�ݦ�񑑍��2b��@_����a�r+CZm�s�U�Ã�є���6����������zk}!���2>���ӀUN�^�͙ݼ6uk������B��Qr�SK��Z�l5���l8kV;�p3۠�ؚY���.��@��;_��x������ET�+_�F��&^�.E�6SEK����3�#�i<���o�&�	L|��2W3�1�_D{˰/�{C�s�B��[����p���<�=I̛��e|̭a�[ڽ�!��ȷ�b���;�a���[��?��,@���;�kI�,%)��W�9~��i�_�
Y�L�885K��ي#|a�0�
���%Co[ �j;�L�:J�$��mX���Q8���ʟ����[��P���u��1�Y �rc��d�}mP2G�7���3)���CM�~J6uc#]���	d��@�5��8
@A-e��z9�s���?�)O�X��zut�)3<�i�Ŝ��Ηa�3���٘V'=�o~�SL���y��[U����{fc|�jMxmD���~�I"1�$_�S{Nd�R��ۮ7��8؟��2:Ͻ���@g���Չ�G-6!&F�J��y�@nA�:�)�<V>o��*u�Ҝ��B�]c�nA��˞.~���	�jDH1F*h�����jv�]�YZ<ғⴷ�\��u�;v��ļ�&���Rm�V̯gdĠP/��[L�sW{�Z/�*3g�W��`����V"ƞ^�K旲������F��l�IMPJ�w��̈́���W|g~����N�(�cB�me�| ��vpDqn+��=���C���$S���r�}��ֆ�c�J� !Ը"����ک������$$!>��@�SJ�c��ң�d<��ĥpL��m�Sk`�Z�:��J�k���n�]P��������*����lั5Vn\�q�^�Z~d����8A;�Ŷ��ix��{biGk�Ab���,x>&f��4�Y*RՅ����x������J�Ŷ��9��Q��=� Џ���tM�����wA~7�1�����o/�1Y����I=��:��v�O�$F�\xˋ���͘zn����Ъ�d���{�|���5�⧹^�R�x$��p��m��K>�\y�x&IW�	JV�������6�u}�VpÅ��"W�����!s�_�1�C�0�!R��k�r
cU�ϒU,q��Sѱ����~����|�����dR��^�۵�K�oUaK=Ht����}�$��w6�@q��Ux'>ƽ��q¬�ӽ�"oBdG��F[��c��������0)(�K,D��{�ǰ�^�u������b��s��(�M�G�d�\����M֝�<&�F9����wd����^�ϸ`$S�8�ҦU�I�N���^�H�`�O�R���;2g}1���}��|�w�m���*e�(���A�/ \2��_cD��$+|�o�d	�Э���@ ���t\{ ��-`	 ��;8bMQ�[ۀ�z���)�w��V���|��}|u����8^�eJ�y��ܟw��u����v��yY���*
�8%n�s�|_{���U��`TD�pZUQU��VD����wZ�k�9*����ހ8i���K+s^��"�A�� 0�
,9�5�����`c���a��/�<i3^!{(�v��6�G�}��c��n,��R��B��;�Ѭl8DQo}�YAjC@��m�6t,e�f����5��V��eM�D��^�^���E?z�g	�@z��6*_���\)s�^K�*�z��?�6�+a��
8�>��;]�������(�4�i�@b��]�䷖x�-?ޡ���<}<���2jab�Q������� �J&@x�lGz�`S�Z?��I�3^2��:���U��F�?jE�lz�^j����ѭ��Ќ� ��2��,k~5>^�,7��� �Z��aG��"AV�Ӊ��|�pE���,�u�]�
? �k��?: �36^1ɽ?�)w�g3$-����]hHR����#;�_> �xx Jg�+.�zn�s�ӎa7��0D�|�� �`��.�a (�  9=Z<Ā�l!�H�S�WwF����a�t|�Ы�z;5��+��-oqCo3EϹ�Bo�6��T�vD�(Tzųɖvx*�<E-�^�S�tor�\�[h%�!m�"���u��y�� �l�-ڭ��ҵ�M�W�g�#@��ֺG|NY |N�N����9t�.\֝�Rt8!�A����7x��#���Y�R�~!_�C�1U]�	P����Z%�!D�[Cɶ~�|t���&�b����X�j��&��	���V��eVS��6}ha��۱@�D0�ݑi 4ʟE1[���Jԙ\�|���$zۯ��筣u`^�ya4���Ʈ��c��h}���p���m���̘�L�nh�_��"|$5z���������������󵹕�1�@�u�L���@`D +7iՖ=����T7|f��`��ęj/��t-7��<�/��m<�3�y���@b���DO~{���g�M��ͮ�L���Qk�J^=�U&�}:2�k�dp���`��8��-�KJ?djc�����m3G7����@.�_�X9d�č�q�l��j��23�"���zc8���y�(��o�� j~�!�ɧ&�j	����5�7�/j{G)�׹�\/wZ���g񯬶
�V,�z�F
�*u�͒�m��/�ت\ y��0�M���j�b~9�2@b���F���� n�04K�u�#�Uo" �F*����UMe��� q.B�C�m�:Cx3��@��[/��,Z��ٟ� ��F�I�� � YyJ$�"`�
Ck2^�(#]]_R��O�p5̛V%D:S�����X�-�c93>W�-,3�;FZ�1��{5YLI:�!� �r����
:MѱÕ�.?D6v��13<�ù HgPFk�}
4�o�	1PW����ǹ��8�'�vd�]&5�4�=~�c�W�"$���&h�����+��+[�Cv���l�t��нXW�ֽϖ�}�j��`3��+�/E��=������P�B��~:�>�Ѽ�{��-���N]���x�0��	�� ?>A&��m��Vk7�(���S��
����j����>v��0��X�$����qU�w�^��?#l��Wn�� Pm@�ۺ��H�%$}���z�tȂ 1ڱY�}l���s��22T�����5�� hô�V�K?n��k9���\����b{9�=��L�X1`����>pe�&��@_O�),e�qw�k�ҸO�Ⓖ�v�57�����]#�Z���9<>9yz��#�O!����j�+�K7�����o��hz����6Igz���Ԕ%�mp�g��Sj t���� �o���5�m;�:}�V)��j�����n0W��t�!�Ȫ���l�z-��y��U��$��`� ��{Pm���[=����*�RF��Z��$��b�Tb����q
�4��Ry�^��&J>�q�7z���/@48B��8����O �(�@0�����Ҳs^KG/ 2�q9��2k\����Ŕ�[~�ó�%	*�s�r�{�u��ά�hMb�a�҉h١�k�-���J��ȟV�ٟ� ,k��&�G�����&�6}C�}fo�0��5�#s�i/�G�����2�f��դ�w�^�O�#xmx�ƛ-|]S�ұ��@�C+��uq��p��PJ3f3�ڎq=V$�Pimf����g7�
�Hm�$)ۗ�T�j#yߒ�����$�/�{U]������M��6�����x@,��ߟ䑨��c�	ڿ����"�[����ﮕ�l~�����:p�G���R�
��E������.�#�b��ꯨkС��@U���b���L҅`p.l���;�<�Q��"�nx3#�kKq���#�C'��7�[�z�s���?�W��Srh��a�GAf�����j����QD% ���Hu	)�%��ӤA�CE������a萘�c`��ټ���g�zV��׳eb�'�#��C�V���%ti�c"8l�w�Us�\)T�W�Lj�e@��8l5�z�>:�O�IP�e5@6֙�ww���$�U������L�C�|x�Đ����q;�E� �B{�O�~-,�g�s����|/e"�S��1B����*eLvD�a���9�4i6�Cʤ�/�j�@vpz>RIa�ޖ���0���.��/���O2|Y�c���B^�w�7{����A_L�"���L��&m������ZMa���	�J�Pb�!���um?R��o�.�����o��9�&��;���Zk�3��g��C֜j��"��@w���b��p�"�*�ST�O��],#��җ��ZI<Ix5��١���7��8w���O�ki�x�!�1K����`G��!	���S�#7>����妢�w��d� pl�����q�HzS�����qdk��=<E/��עBg��S�k��:�dk	����'Q|�Ou:�{���ݑ��˳1:�#Mx�0�����󹤭��s]$ޯ��-����bI�ϗ*Bax��IKBP�P��w��7!�2�s���ե��ѷ��_&��T�v��ՍC����7��"$�g�QW N�ON#|)۠x^���9L@����ό�9��>=�~���"�&2j�E��͗c��=;G� }䫩��:H�u�M��������w�:����9�G�DŴ�zS��M��8 �
d�
�W�� ���L�u��p2��8k�V�Ua���� E��o��������]-/(_ �;*f�:�x���$1����>E��J���D*�C�4��� *�_(�a.ں	�_��<2=/�4Ȕнt7'���q+���R��T�L��+��>�f���K@WS}+&�,���r'�Ջ.�ڭ-j���対]�x \�M��om��/�?tD��Ҵ�a�T2������G��F�����aC��������9�������<�����|��C������~�WW�*���63���W��jFR���T�[!�}��0�`� ����p���=�W:�M�j��V�J))>�x�s�������ѕ����8)/H�� Kc�����ξH������bR���#.Gui����x��"�/��)�����q����U��6���]XFo���CP���f"��~��=���щ��e�so�"J= )�Yq��n�'&��C��������/U�8�������ѷM����]��b;y��K{���D�4�l1��z�5U@â?>�t�$�!�Z"��毖��u�s�o�Ju!� `\.��X3@��e'y�姀�6�C�@���\��kL���ր̃V��].&���d��{��kꘗ��1<11Jk@3��|�ƌXK�%̊ڪ�.ꈺV��>'�eFn��=���$A���T��c�:㰜���=�֭Qp��i'C����l�]BRcQ6
��v�J&��k�YΛ�������!	|�@�9��X��4Kį���@�����s�����- �d��d(�0\ȕ}bc3�+��z{/��#���.�o_�:_a6H�WY1���"V�����$��gD�g�pݥ��O��`��6?��$hթ���w��Ϫ'$ߡë��q.=���Y�k��l�g.RG^�EN��n;䀍W�K$�(�IUg)}"�'@5Aq"ȍi�ٴ4�bU�X��������E,�F��j��,���J�}q��gM:�Q���U�_��;�h��pՂ�r��~��;�t�I��J��z����x@,�Xsn�I�0G�7�1!�H�]�%z#��
2e�!Y�W�Y,$Iy����7.��Pb�R��Fmjq�UۺmVmH��t��k4����6�� [�0~��][�758x+^���U�9_H,�;5'E]w��㙘�p��ԇ���ۍs�� ��n����5��N�J���ԟ���7M�u����z���~\@�+��')�^��^�/��P�6��J$a/��ҺGآ�c`�a�6���#�m�E���k�_g���u��=;��~7�#�
�b ��JR{;nNf6
L"&u��@H�E��`���
/qHLQ�
3iZ�C��P9�\J��d�vK�GE�oes�k�Ĝ��NGωB�D�נl.d�=�����?�e�����= �^���O�V�d�7�:�I���oU�|eo�̮4�\��|�U�w��'���_4u��ؓO��E�;=��~M	q RA���?�'=�!���`�S��wR��bM���\F�G%���X�yxYp��Ӓ�I�xU�Z
�\^����Z��Q�5���'8��hh�����J��0�^oڲ��$�y����hrK����^���e��ྮ���M	t��.�PA�RjY�[/�־�̜.���;H4-g)�`v�b��YP���L0�����ĳ�[���&,��1s_��]��Uo�s�@ۦ�f
�ߩ�g� jQ,����j����Jsԕr�7��< �1�����4�(�.�Z������lj	=���\X�[]�)��T^�H�L'c�?�|6Il+c�`(��x`ò�����	�����F|J跐��p�j��x��A%<_�e���CE����;)`Pv���#4PZ��������c5��y�V4R"����Iq��饎���#������;V� �0��!u�^`E�r|*M�moc}�ը5�?@���g����'V��� �ʽ�mm�E6fe�r�S ��2-�d�oަD�.�6�~�R0�,�F�
��eq�0IK�b���V�������y��:�p���3��|�Q
`���c��6]�t�k�W�\�W%��A����B�3�+{r�E傧�������P���o\ QD^��3ɭ��ݘe��9 �(VOH�vބ�l�J'�6��������Q�Qs}�R �c|��6ю���N#�U�>�V���P���k�G�r�◻���K�M��`����ڳ#� ����mx=��sQ�j���?΄�7��hu�.�A&Z�=�K�j;73&N�T*�:�4{�̖�~;�_Bq������ò��a*��審X�DA��N��Ԃp�G��8���@���fX	�f)���!�3��p:��9��[,��!�JW��xpq����ǉ2�ne��an����1�>Y�ܓ~k_�ɹ�C�D�@o����*��.�5ww�q��
CZS�i݋������l��'�PP�1�i]l�C/T��.0�4a��"��>E�Җvs�ƺ�|���_}S�3���X�݁7���Z���x����֩�dU;n(����%�<�p�T!>y��f*<�gO�О��3ßkMz�;:A���{�ۓ��{^NuF3��gluN�%_�e��F���߆�W<������v��1�M�1�>��k�ts1�3U�M����ZP)X���,�:`y��i�����U�q�U�M��a�����4��G��J���ӌW��]��y� �.o���m6�D�G��"�n�^mX|�_�Z�5�x�ރ)���w �[��5��~�rs<K� �����}ÏzZ�΋�Ğ���kkd4���*~��?�[��9%��j��������5�٪RK F3g�B;�p������.WRj١�JNƨwŗ<6Y�IS�{�D��J	{�A�����/ډoW�hbc�O���Ԫ���ݦ�;jRJ�� �Ei����5�]��!�{�s�ݚ��
a��W�,~��6��ԇ_�l�?��_2-��pou� ͼ�.����W�R?�v�gw�~&�&�}<���:��#�p(��\*�!`ۊ��c;�c�\�6"�-^��`���}e/��`��s+�-���O���ձ��`�~����;ѕ�/�5�@�s�Z��q�8y����<`�G���b!��'n�MB�w�ٺ�q��^!�ZS*ɋ�����f�J���Y:��w�&Y�Ք���>�p:�|���Iמ�5����m{����H�t���a59�.(,���|p��7	�F��$�%L*�xw?�x�0��V�B,qݺ��BIJ��#�:I<�xi���M�pR�v�������Z��3�Pn��m�rlt���6�'�|����TAv�܇J3�W]f&?<���틧������y�Mhz�O�P�궡��gW�����5��3���@±��A���o6�6��)�H^�t��m�v�Mk�4�W	��U�qDJ��TE��k^�m����d@��*�RMS�t�|�C��!
,5���� �"����uPt�/?�"�;�G*'^&�X?���Uv���n��J�9 �W�dui��Ο����o�7$M��Y�ʤ���j����{9 ��*�܍�uYA��}��f�e>��g{�A���,�L�AR��z4)6p��W��_@g���u&�]p8$�|K�c1~�#���&"�؀p���J�,��nQa�Z,��~�:gZR���|�~5Y�c֥�[�"L ����fpRyW�l1�a�0�,ITB�]`��1�|���e�y>��d���qw\{�F�?��]u�s2t+�����AQ������j�C����O�����M�7f_�Cfa��d��M��E�%l�-����(���{���Д�~($R� �|/޹ы7d�	<�:�~p�~��e�>{4�ָ]=	���0�`�p/�k``i��w�Vd{w�쎨5!�7�q�4�W����$�]��p��Iv�&��0,#f��0���\�!W�q�O�_ϳ�%��>� �xP�����,e3x�Y���~�JQ��5?]u�B�c9�5�������W��))�J�qڹ�?X4�gX��F�Mk;K�U���?[�+D�o�R�jZ��Y���+�����������BJ#�'\SS.+��ύ�4i,��b�\�B�$'	f���5^�p�H�[6��#q��i@�h�݉`���;�N�U�h��%����'��S��k�'I�ѹ#�����9E��zT�E�u��1U�L���v哅k�
�$޲���қ�)<�b������ScR��q�W<�
��|���$�������vGJ��/�lU`�<o��
 �l��ζ���']���hh+.�'��Fm��&Ɣ
���ʟ��L!hZub������v�K���f�'QAb����5��7Ԝ@�?b��+��?�_~����F�AZa���b|������:I�9e������曏��0q�ߤLy�P����YT��a�Y>qeZ*�=�I��Ƞ9������Q�@�.�2�Q4}Dt*�����zc��j��X�@j?m.ȏ�)���E��"c ݦ����'�P
 �J)nD��a�'��L&;����j��m��p����T��<JtI�}_QU���l�0�}D� ��!��>�� zܴ���hX&��i����v)�rן�V@��t�|n5��vk6�M���]���אں\"����˚�"Lݍ�L0m���������=/E�\�ܖ?�3�?w�:���%}�5�R�L�oR!�3��<X�����a8�5�=���q�����Xm���(<h9ͤm���d��''u�
?Zw�
D����n��j����-�� ��}i� �u*ӵ�����<���;�a+ҋ���昴�	 �D@仓ؙ?�F�#��7Mq<N��Н*����y�+��R��X�Qv��c��R���k9�`/�G
�G6�D�2"�NZ��D�D�5T%�6��қ��A��x��x��vv��p���"7�
��{I���g��vo�q+�6/���T���Fs{�;VG� ���v��ݿ(��,`U[�a¿j!��X�y��$aݼqCej������������������eq�᧸����R�>�$.�&$Sw!�W���v���]�g:W9��]�;6{�Y5��������c����Cfk���Q���ɜ4�VKX h���F���3LT�d+̼���u��O:�~<�[�\d*ڹlRؘ'N�$��j�xv��r<��.�x��W�W�+o�2~6�U�"�Q���@��V�-:��-P
�ծ�����w!�{�=��ߢ +���	a�y���.�u� Nn���`�CQ2�@�����PR�=��h�u��oq���=�·��}�ڌ*����.�8�3'�Us ?1}]%ַ�UD���&	�������Z�7����0�Y��p���.�� ��$�v�zZ�3K�	�4�q�vF͘�R)���6����t���A����D �����m�^Q9x��Zr��<$���.�m�{�hbw�f|Fi'8k��l�7�����T��HZD2�v�y���K���a�D'�O�}+�d-e��N55πO^�T�9�.�u��C��Ȓ(6{��ߖr��y����X*(���o�ʣ&��`���hK�A�a8�����9ňC%�Y�#�%~��,^����H�K���󂖕���=U�2�����f�&;o\O)�
\��V�����l�Rm�D��i*����_�dn�O/M�NHDy�ރ�g�ʪ_1��~�{ŗ���D�,<���ހp7�~������b�ѥ&ƿ:�^K�;��;I���GL�)���;��l2 �>h	��^<�_�Ǌ?��<�nv?8�h�	 ��)�ܳ;I���t�Ip8��n2��l��K5��c�M��l��r:��$�����/<:lͩ��:��3?���	�+�1I#�q�+OZyh,���|�2*f��B4&S����U+A3�������#&��K��!I;-2��Xk/Y�?��,,c<~��P��N�����g�Jߋ�W�� _�۪����0�^���������s{2ԉ�6��Yx�B���u�3������U�>��")^����߻P6v�w�(�gq�����;٢閖�+U�g��0�6�`%n�b��� �BS�pIд/T��	0��q�Eq,O�6�P�����2��Ŷ�4�ڸ���F��o
?�xgąT���jT�l7���M�8|hZ��cw�
nw�$ou6�w����>΋ �g!���?uU�&k�f�6Z��n-�s_�MOƃ��_Q}���Ԇ_q�2���M���c0KT/t���9�J����ܨ� n�� Wqt�$C�Ѻ��@�ä�T��ەRf	�����R�����Ei=����䡥�Kx[Q면Y`�쨬"��*L|k۔��N��۹p�}̬^�$5�1��}`��>��5u���K�`�j�+���;���S��} ��N�V5�]���7F%jNX&��Ǟx�����.�v���lX�c���:=���J�ܧ����4A7��S�*"��YHd� /�j@9��Ϧ~g�M��2�j���Ϯ�Z�\��ܚ�\�Aq��bP*A��n�e���$�mQ���߱^N����JR}\Ld	"�-�yr���,�+5c����ch�~�@ �n�'����o!s���v�����ȯd_���������na��� #��;M��;����o>����e^��sd�A�Ұ�!�|�o�_���Tßr�7��Mʝ��
KgJo#A����}}3v�u�OF�J7�����M���� ��`�ΩR@⹧��e�b��^��F?��jL�7��D��S?B�m��Vq|�K_L=������`Y�x����2r�q�l�:��-<d3�Ld��J���o?0�5I��	~�o)����YfL���.A8��(�w��s�x`��nmx�����x�����{��m�k�K�L�1���խ�f��M���ժ���H�*�ݩ���uV��8:��F�!�Ӭ<)*���K���4n��o@{��dԎ���I�3��|-[?��� �����Oٚ���^�>b;�c`j�yW�!߭#�aL��i˔�k��jW'v���S�X�B��SP��"�ͳ]��y*�p��Yڐeè���
�AfN���
�����[�>tZP���~W���i�
~��~�4�CG�����N�ܸ��mg`����>y8v��K%{S��ik��$p��%��W�5����������A�d�LĚX�y�g�?܋�������c���c:'�a;�6]�(ŗd�?�L+�&����^�����8?���=�W��zyJ����T�w���k���P0a-{-�Vm����hU�Um�ohjqF� �Y{�Y���y(����0Nۦ��Oϼq|���+ǥ�O���o�UӔ�8�J�����"�'��8����� �����;θ˃Ѳ���]E�}���#g����&*I��7�a�	%���c?��/����S.گ^L�hę"YhY�oܔ�2����g�F��0L�LX���ag���������t�Q��t�f�m;�j�˷W�x`�W��P4"oc����~��CT'-M�`Y�Ф���7�O�ߝzA��i�����!|�����'?v�lؙ��dr�D�"���t
�;G��QċW��Q�s���_M1�x�P�ӿ�S?��b�x��z�qzm�ӣ�PfR�J��$�a����~S��E��L�Z��M���n�E�s���l�G5���)����DuHm�J@B����:N^�Pޘ"���>8f	�F�������oM��\c��	�.�Ac�f��G��m�l�吤H���X����ܼkpU'��1����ze&��{
�����w�@�/��wa��t�`��>+����Z'���`U��m����f/���D�u�"�Z��s�*p~�ϱ��/"Y���ސi���u�
A�-��u��;�'����ad��˯>��P�!���J�}ۀ��$Y_�m��k6)�-�Aua,5=26�*��A�����ĥ���>�a��Ǎ��E�+�u��l6�M���i� c#�F
:iI������Ք���hzN ��1	���9��!"���2�_�����H�c`�iM0{�7��Ja����?s��+M�m��@�S���vߘb��)��	Aggt. 5�WX�@?Y7�~��KH,�zd*KZ|�x��|O��p������cM%7sN�)��9�sϗaA�K���)��y���7�H��%9e�e�	�lL�ǳ��S�F��sළ��h}���k �ܹ���_�^�+�e@)�(K�8�1�������^\�]��U�m���F�w�d�|B��M�0��D�����(}c$11%^Y����WWc��a\֡��RҽM�J�!�m'����{��Q2�XWW���`���ف[���ON�Z'�8�*W5�L0�d���tq>���o@�@��fff�I��p���!o�3�
*ۍ��)A}X���b����,_���~Cݛ����ܤ�r��/�o�@j5���lJ,���zG�n����.T���r����0�G���F�Lmޜ���f'�u�u?<�h[L�O��8
����\{�p�t50��K/�w��D��� L�'�OA�� \��o�6�'�#��ͽ�P^��]����ng����U�r�z�c@������`�O��j
�`�?_RW�ʼ#���5z��y ��H�O�$����b��_D+'_��	����)	'@0�IAh%����B!���� �7�$R��rԕ
*Pob�ݡR�� �|�fl�=�.(��x��r�C�d]�0:a�::��/���i��H�is��s#'�AM�E�Ӛ?����4e���[���HF��#C���
�s���A񤈏^ϲ;�u��̊���t��6�~T�
W}��	�O�N����M�s�6e�R�1Px��
�x	��a��$�x"��e� @#Y�*(N�昷iZP���l��v�u�[���ȖN�Z�'�ꕼ�xd_���n�;	���uQ	L�Qd���^����nu��W.�*7�w���S��Z��Nw�qA�e��q����R�d�w�OJ�;�Q� � �{��ii�
2!�Z�%�az!X��KH���a�~l��+T�׻�_��G`�#�4�"H'1��S�;Q_):Si�u��V��c�NY:g��\̫��ܰt�k���ݔ#0��@7�o]�ى�s��b���U�Wy^�|��mN�����;��o���Wk<���@w��/(ߛO"�W[���,��$��񱉣��	@}�-H���O��u}Z�"0�+[��v��m���1}�Z_ҁ���w(:ƈ�4�G��eGx�.1X�p�a��c96՞��[���Q�U��׬\Xu��H��>����J�P������gҠǘ� 6x�Q�j���=Kpz�����@�bY��'@���++�N�`��b}T�� �_S])�<��7���$@�d��޸g��}���q�I��JQ@���_�hm�f8 ����)������p��8����*G}l*^o��g[���0���\�6����j�A~�S�DmFQ#W��P���r{s0��%�������h�ԶiXD�-ۘ��ٟ� �� ���'&E]2I?���Z�fF�T%Gٹ�{�[��r�r�%��Bn�#�u�[�A���Eg�۴�Y�{�4l��X�]��~Զ�W<��bj���V��˯��!����<�\�['}S2�q��d�� 	�����DW7n��p1ֳ��80lCC�>����	��Y��X�/"V ĿuV��_Ⱦ6C��Y�4�}މK��՛���I����̡�ܠ�xL^g*�x��叔!�WRNۿ�h��By�T[�s�B:�t �������?���5^Y�)�c>��fi{X'��ҋ�=m�DӖ��;GưT���3�0UW���q���h���:�}�tr���L:@&�S��� 4@g(]�E��'��r���.�)ծ}�sJ+}: GPVnQ�v�$���I������!�ޝ���qȝ����r��ގ����µ�Zm|�a��9��f#k��5���rW�lu�<^w��h�j�U6&��2�%�<�����椖�>��8�Z�7�N6��6zX��_����$�'W�9����!h�9=�0_���|ܰdh�ȫ��Zk��죬��d^�\�|�m�`�O�Z\����<��v9?Lr;��_��E]�M��U���}�;U�>�Lpn2$��~Vnh�`b������/�2��� =W��!粦f/��$�����u石|nwVƛ�=C&L��^��₅�x�-4���뿄gz�u��m���v^�Z�4��)+�����Uv�}v�l���֣��T�9��&R-]$'m{�0��mW�Y&0��QB5Y���C�^Ub�.���d&�Vg�tE&!Ӊ�L1�
ۣn��H����N�[�D��>){��+Ob|Kv�Vu_{<����S�a��M�������Ґ��qe��OV�u@�<���2�r6e�x;p��˳s>�h����8|�f��Y3�r1*Mr?k]�dZ0b��@,�^*[����[�(!�^��>N����:fH�H�����$��iK�>�"꣥ �g�p���٣3���5K<\la���!2�x��l�4~@Ur�]T6����F�����&(�|/�r;QA9{ 
�:G³��lT�u��%��Z^�S�i���ai��&�2A�~@_��A1gKd��6�[���/�m��>�L]�/�ds�փW�vS�QC[��L)��p��	$�$�P|nH��4�H+AGX᳒Z������L�S�����褣�>���N�ቼ���n��L�W�O(��Lu@��6���䗙bZ�њ������ϥ:~Ya��E����˃.ee2����}����K��2��yJ�m�:	>�_���7�<=z����zz�Đ�K�V�j����ۻ:t�Y���zT������fg�-���:@!]����)A�����k�1E�"˕^e��ύN�Z����g�x����t�h�]t��&r*YcK��`b���m��saIA����8��%X�GDk4���I T����>���J=#��}9�_�/3�Yhx-�Z�WL8t�,?�[\�:�Ջ�m��-W�e5n��z����j���3���堞��[T��r)j�d����Az={]5C7u�»O%KS2!�S�����48�p�c�M�ǳ��
m�hM���eR&ݸ�I3$��!���w&�#�?T05-h�ط�Hg0G�,����E<�^�"�l�}Wx`��J�I�Sɡ$*T`��/��}K0���j�`߮�J�q��?l�I��,y����v���[y�����S����rj!jA:Q�S���Lf&�o	<�c�7�!�y�+����6-�	���oۍ+,=Y��Ҳ����ziU� �Ʌ}A�H'5��~1�^�"� 
{���^=�0�n6ڷ+vs������s�+�g���1��K@�'���l.������8: N����ESQ�[�
�:N&$���e�s9�o��`� ˄��a����P������e�MN��UK�ȩN""`i��(�,��@�Ȫsn�x�Rʄ�{ҿ�5�6��R��:����䀠W���l>��x�B�ۛ�Eݦ�=p�5~�&j(��o?���B�962��Hq��ۊ�G�K�7\�o�����W����L2Br$牟nnf�Tڣ0��g�y��I�f�!���S>��4��I�-RC|�S�u6nMz"~+�;�B�mh�oS����5�b~�i�Wr�Q��l�D>ǈ"Q`A'�.e�%y˻C�G��#��hݳ�_ah}���O�5e�C�ZG?�����/��.��+�IYv�Cv�L�~�4�n��hO��*x��������,TƘv���8�9���@�8���\�<��,;��HYsF'�-��8��aVT}rIu[+6Dy�~Z�]�[���a��h43�Q�v�-@!Ҽ6&>l_���b�@�˱�QT����]���5��2���1]�̡�fZ��d�3G1c�IE7PIt�ы���*0���N����"�,u���5��K��c��^t�U�@�Fֱ��y1?�R3W*�����ƤFg\��Sbki�+����K3����I�a�V�����kcr')7^^^�y�9�Ob��E��Lg�}N�8�t"1�ձϬ8�7�=��+�~��u_����n��"i�-�[��롩'�2��VCU��)�H��x��<M�ը�D�.��p>=����/�&��v��>�E�d&���Ug�38U�*��!�Yw����nrlV:�e�&��M�N�����M�]9.�Q�Z�& Zeq�����I��n�Ȳ��Ɗr��pb|����5����2~_Èف����	py��+���ݞ.��~�X볃X��6Ƀߞ��,m�o/�(M6w˸'���Q��N��µ�T��(�&Ɠ�"�)�,s4���\ҷ)u�0ik�L��Z�}�?'f~&h�=��u?ҴS
��~
��a������[���py�U���Cqz�$�<htK�p�}��@<UX� �,\;cj���*x��GL�����'�r�DM�=~���{�:z��,08�����[�� �{!�o|�H����ZK$G�%��x7T��}�C[��äo���R��iP��Jd��Mю6{�9�ZO�~@�X��|�[W�i��=^\U|��&����o	�p(b��۱%f����.H��M��Uk�5�}�ZG����+��IdVN�CeL���h�<�`�*>0~����T�rSbO�"�ҩ�k�M��Ob��jk���&��ɑф�usO����1PJ'	2�:�D4��[�S'�6���ŝF�=V�=��:N������o����y�n�b��qߗӽ�������Z��:��F��/{N�M�ɗ35k�$QyZ7��Y�<��n��p��44:���:��{+�W��<�#�z(�e��`�|U_�o�e�����X&1�<�p��.��/���{c#��E�~u��;\:e���D���b�(;6����eA��\��[c��UoR�F�<]İ[A�3�|^~�4�z����(8�Z½�q�\�l!�����}����۔��ZU{(����왻�J*���|�)�o���m��#1;,��X��~���j�C��	��^j������}�w)�T�Ͼ+�����ڛ$�϶ě�a�G�_��&��u��.��� 4-U�8zU����#�'�9��b�Nz>]x����{���;�)��Vy�tߝǾ���8RW��6&�գt����Q/�԰�U�<�ZV��%j�����>�s�������D}��zie���[�T�n�
����y���2��)�����\`�.�w��J��+5���=�Z��tǽ�u�NQ]�����S��e?�p����)c��ř�[����.�� Ӎ����E��_�18Fs�y�R�,�� KצU-3ӣ0�UD3��L��Yʺ�즬�3�9m����u_�Dl�ˌ-�,��W�P��/�&l<j�7�*�C���Ḩ��Խ{�Lw��S:(��ט*{+ ��O�?7+F�t�t��ƺ�F�7[�n�B�m���<�����3�%����訨A���嶍��1�v#U�Z8���	C�2d��Pj�ͳJ���I��3?��M�7�dD�p��/)���������O���w�j��Օ�����7�*ta��A����Fle��k2E�p��R%�PpOR!�V���*m��n;u�Uʸر�xs�͛�_�U9C~v"���O�T�$J�҇ݏ�?��6�4J��+[�#,mK��U���ޚR�~Fqe�k�������|��q�c���:�0&�qk�uA�Ã���#��2Zw��&牻�E�z�H�1aldj Kʲs�~⏣�~�}O�M�W>�s�j����g�wa�Qf"�7��ԆY����^���D?T�Rm�;�qX�W0�6	��%���ݹz����y�:���a��������$.��%���*��ȟ�j{�:OV-M���e
���7q�'N��Wͅ�ll�n�Te��9IE�*�a}k,�\�N[7f�E�fy�xO�類��=@�-N��L)���fJ#�S@�Ӯ�ZW���p��uٹg��m�k 6����;���>)�������ʔ�[��lXWTp�,#�xm�L��)�:\�.Kl����f8 7Oْ,��4D,o��?��u{��{y�Ξ��]џ�����2j�5�o�N�����*rm�XRo�ŝ}�]�Q�}��5�`2���~*�߾V���ѝh
��� ��T��
��6�!c�,��g�;�f�s#���n�j��{ޘIkv9�8�3�ōo��˱�T-�:
��2����A_�K=͋����!���;M�V�;qW ��ߪ����DH�U*���#V�ٰ�E�=BA�pc��Y������p��u����MiM�++3��m�m�����'	%.�4Uf�>�Ņ6����R��%zP�|�^# ��DW���S
w?p����h�E:��P�b��稾t��1>ŧ���݌`޽���3��LE�/v-[�����J�$_��Y��X����}�1М^�9C�M4g�]hJgTՙ�x�xb���gUs�Z�nS�K�e��/������1fJ��X�Z;U�r�?�hP[t��½�>]�����#`n;�s����N��c��~����!-�ISwף)oܢ븖��J�O�CS��/f�JF��jd��N*��?�VN���"ꃫl����3��O,#3�Z���/8����>���g�(�=�����ӌ�ޢ!9Y%Uj4���-q���n��=q����[=��rPA��C�6ϫ��X���f��1n2��1��K	z���Gڧ��"I��8|����*5?�r���j�-�9�oN�m�Nzk ���>ə3�N/["��m�n{��Y����kB���з���M�4��u-���v���w������X�-��^��gU9r2m��J��I��u�F˹o�_��fkG:֘hw�?��}_'xkk�=�Z敆�㝻��v�^�6��������/���٥�L����m�Ԉ-��w�e%wߢPߕY,S��s9Yg0O�F��z��Ú��]���d�:j�AK'3�)i<��I�>��is�[�>���JU����:���	-bJJÏ���2V�4�$W�1��J�gCݓ�;��S�#!��@춸s��Uݖ���]��J>�&�s�P	��u)�
��޴z䅂���/9E_��HH��������_eV�:x�U���c��,`�}{�2�zpq�Fs���94P\���ל�6�+�m7�p�b~����HG7R�3�^��B���4�b�B$�by�?rAc[چH����\ק��'��^oV9��7j"���¯(���[�#�{�=�c.S���2y�_������ݕq
�oH�a�z�
�����I��x������:�~��~<�R0��:�
�e���ܶ�8�m�و��Z�xL�3�_��W�i��N�Jޅ��xP`��Ʈ�ɥ?�FGm��Q�߸�l�
��Z~z�ހ|�R�)˓��k')���#��Ȕ�,a4A��.�-�y=7�3�=B�%�5�(C;S��P���/�c�'J����gݷ��+���BO��G<49i �O�Tb�����6ƙy�_�'S�����ɧm��a͖�нE@�Jc�I�v@>
�ngZ>3�+�e=����Ѵ���+�DR�>E�xDN.�K��`y^�x���
�n�D\�t,����2��^D++}��NO�����+锋B";�Q���~v���&�櫫��=Z����g,Weo��CshC�o�y���M�R��om#�eO�B���w�V�ٗڱ�+�x�������H_�|��%´< � lW����#��O+d8⬘:����a��ct�O�	�e:��fñ����3����A?E���b��)����P��m[G��J��v83�$�^i��C\b簚,�T�Ы����v��ViP�mF�����vw�t~N�K�h'�m] 6l��!��
���g������#�� ?S���/��� �N��t2��L]���LŴ�m%��&�P�|��ڷ[��6�9��:)�Hp:IH����R����?�������k�7�!�a��Ώ�@��cH�.�^�H:��G�W@U�}_�	�@Z�)��$$	A�C:E	)�CB��n�HJ# �%!q���o�{��c|w�7��}�^{���k��}G�R
E�G����k���Ն{�i��	�r��޼H����3V�Z�n��y�V�q�>���6�����ZH�bhA��y�{��m��ٍ��N�hl�7�A�)�h$���
X���Z�%�6���� ��m�s����怦�n�2�ÕZ��-2�$�����?S\��V��J |C�L�7��%�:|�*�oU�	�B��&ҽ]��HS<������2���@������3��Xj[�#t���f���z៬�GL�{Z�WsG���n���� ��ʯo�F�p��
8���]8�oY�������v�R[�S+q�pR��>f7f3��[��ʷ@-Y��o{�{�����0�Z��
���cqgQ��(y#H��b)�g8��x�t�@�t�d�=�cf	�?��.i���Pc��4��2��u��?߮�D۞�j�S<|�O8�`{q��9#�����
ZU�-ֹ%�8�D0��HN7�|"A���(g�K���@�%�vZ��h���'
��>	'�p�V�*N�jv��w�A���ݱ��}?�F�i�U����ѷ�D��1�&O����϶�5��ΆtDo�IB�/�4%�k����w�[��䌊�nlÃ-N>��I��F&V�I�o٥�S�n�1H��\YϺ�4>�����̝��q�:�uLN5��'�1q����/���U2���
�g$�Bn���L�6L�-L����`��ڽ�	��p�M��G��=��ñ�!��	>�w��G���*����RE�
������W]�a-�x��wXr��b���-ajp/
L��(��m(h��W�&b0[�ľ�6x�3��:SS6�����?�ꆖE��;����#7$�\TJ�+���ig��,��]ߐ�{�9|���qkR}�ȍVN�J!Bg��N!�Y;��x_G��p�9 d,%�-� ��EUt�-�1�1u7���xj�W��!��~�e�)].�\�#>k��B��6��87���П�c������o�:��wy~�:�%=��:��w�L[�?������`�é�����v~�j(�A�J��k=��:������i�9� >toU�����/=g������Ѣ�j8Wg���c����֫i�W���� �^@B�fD&Ji����
�[E��~��~s7��C�!�488��%^� �s���v���Kw��.������@.o���1�Hq��	�9��m��|�����٫�r��;)�@>h�"��I�43Ӳ� nɏ���v����]��\�(v�*��߿���'�7=HFnؼ���}��<��	x 5�������`������Z���9�LΜ �)qn�U�?��}'nL�@�����h3� � �7|Vk}�Zm!"��e��n��m\k"7/R
T:rjc]@�,M�m�K���o��{�Ƿi�U�t�S�~�s��즼t_p�3n��c�?��%��ܴ-� ��/��;]#�$�\$�qT�o"L���W#�1A���'�6Fh"�C��ʹw&�f	C���[��K�KqJ9��3?��q�zB{����G�F���~ޑN���ڛ(����J���7���-��D��}���1�`F ���t��0Z
_��1���>�6;��8������pc�ڸ��
nzq�]��ǩ�6�+?�E���힆�"�/W� h�Ҷs0_��v����.�@�*��?�2H�y���������[�ʌ��#.R~ߪ;�}wL�m���а:�ЏO{-�X�q��R�
�7F���٧s3���ſ�&D�M��v%� N���M��DG����Ȱ_�V��8�#\�:�W i�o�t����QM��to�,!ƭ�0@Dk�|��ƿ�aSl2s�A�����<"�w}j��@��ڒ��k�t�&s��J��DB}l�al�괲��<G�oCr!_�0�_Ť��-Xn�� \Ap�t��j��A�#R.��Q%��1�hŪ8��E�$�����j�M��a�}%��:���e�Ϙ�C��Zn&s�mⓔ�Xwǲy��j@|�ݨ''�����R���k>R'͸^PgN���א�Ƚ�'	�&X�LO#�Ú��[��i���s^j��0P��f���U���G�#������o���%���u��42���_}\�J6V��7�M_o�#=�?���~=MM�مk#4(�F�Gq��JI�p<�w����2�[K�;�R��h6(�fNx�`gd�2���,�k٫Z����¼���Jo�v� к�TA#]8��m�#ϛ�չ6�/B��;t���1���;�
H�AGDY&��d���FS2d�;����p�
��T��1#�;��̫�~n�+�\�<y*����j�=v>u+��/��U(�!�,1}�ýl�W�v�"0�\>����g>�����C
_�!7KM3A>�0[����0{)���`���p�Xz�!
��,�V/��KMg�#=[��)�J�t�'��Em�Iq0���Ý�:'�����qQ@Y��YaQM����m��^a`�5>�C�Uq9�2e�x�':a¬�̄�S�h��v6�U���]�
����\���4Hs,��B��V|��U17��G_f
_1�~��e�.�-������1�i���g�iQ�G|�?VD<��'1K?�y�!}>4�����9'pL���H��&���R�:�Ua�y�_�(�dM&AnxBt��T�ϡ����$�p�� K�)��?D��ϫx��?�y}�9W��'����/S/.S}����p�ET��;�(t���t�)��q� qA�s���f#��_���V�RN�V8�H�4�{�� N=s�X�֖�i��'����w�di���#٦g����ʳ&�l����ˡj^?Gi�$�A�a�N�g|�ux/��Ÿ�E�!_z���% ����̄�%(c�ǳ7���l'(9Ll�3P_Ɏ�L����͆?%���4tC%�Ø�b�M���I�fkd�����7_�w���W1�e �7�:-|���d���R��'��iD�KB��f�A���ql�_7�T������1�H�ɑt�1��K6���H̛^��W�K����\�?��
H7�[����J@u�-��/�hoQ�|E���:j��#2;�����X�����7�TA/G6Q�R$S�\a���� �u���94�v5��ذ?Ip;_�D��1�+,��")�N^!+�Dw%`��:���sg�@0@��҈߯�D �X1��E��?��C`�X��i�xJPR8����Y\�؛TLS�k$>�/,}L�Ql�F=Й�">�-蹊'�p�K2��^�{ b�V{~y�|��^��+��J-��]��~h�

SE^R�х3y���O�Jƶ��ߥ�2)�}�Yr��9�H��AQĞu۽<�3Q�69��	|��E1f����*I!R�G&�pÛ�eK9L��͢�5ΥY���&(c��-�/��{�;�~y��uἹ{�����O���������r(Z��kgϩ�<��\M���U������G_�x�W�g]�/��~��Q���d7���Sg/KWvb��v��?+�F,�G�n�Ir.���{c	��<Ț�
q�޽o-����`�!�#XE�|�TH~���ջ0�7U���;�"��s*�����=��zRVot�T2�&:;h�B�X�����֋�`]�4i�5�4��v�Og�BX��tX�r�d"o�
%/�p�P�Y�Q�WLʋߍ�<'�.��4�r\F�T�YfJ#�o�ƞ�����V��)N��^).�}P}kCW�S�ۭ� ���ø��~Rd�<�|��<-�ӫ������e?#ۻ�z%\�t�5��Q�^�������4����#�&��qK�3_s��{{��B���%j�����ѭ/��yV�I>����2J�bI�?����f���	m,�%���Ν4���?�,�}k���v����+O���A{�_�y|���R��m�=Z�mn���5ۢKa��-j��+�S�@�����6�xj��ZT�y�^2��̈́�e����#���u��i�0����]�q��svm���kJQ|&{Go�U���.xo�eڽ^K�jb�|k �aX-���_*O�>���w�i$�!�������F�v]c(�7r�j����@l�a*�讟?m������-  W૵J�t.>�yw���]�~�"�ȕ�W3���)mKZ���UAz�ߟ�j*�E	�ˢ#׆����lP��ķؗ�뾖,�?��*�3\�bi�Ԥ�!�__��F����"�"�2��M�rB:>,�p���XS��>ڱ
:ވ�U$����:%r�ʲ��kf(����,]~
P������T�B,�N5>�4w�y�2�3U���j��K���n�i���!ыX�*�ݏ����"�8�R�����+i��v
X��>�-�M���AF�sm�����n���>�(WYr�:���H�KqJ�Y��WL�B�\�u4mL�j��W�^�W���t4�I��9W*B�M��h[P�J����@@f�*vNyJ��h��;�#_N���fi�i��q:W��bE�����)�Y���A͏���=P�2�����DMN��1e��ɥ��O�K����/���=Cs���A�#�Dk+�������v����~y��{� ���}w����������}���B�4�i0��e��M]����E��^�y{�7��kz#��˜�/���w{x����dE��VX����q\���J��=�]�E���G�\�$.��� ������������|3+%W�U.`0Ҥ{w��*\��=,R7>b��+�
�����3��k=^�Bu�#�݈:Jut4O#�����mi,.۾��z%f���W�^�Bp{�
±��X�������^o/)��ɖ��Q����Z���T�����.ե�?`ZP�B~����Oݩ�99���Ͷ?��ֻ)T�Dؽx�P�U2$a漨�Ǽ��b�͋û����.xû7���0���������VC��7�Z/�婅��[з9�/K�ݽ}��<u�� �}��.1��	�9�Ѓ��][�&�ٰN������������ו���<���׽2�4��6!����8��6�3�h'���+A�����2!��>ՠt:>5~Ԣ���;��_�u�(�~\~}#8���o�lA�{��K���gh�m�x�/faں���������mN>쓍4�ĘW8_��p�'�O����s����a I���d����z(7m���S�U@��ޣ[��
�$��:B����Y�����e��%���_!��.�LR�@�G��^�PF&�m�!L��jb�����5P_X�'Q� �K�n���΁ �Fs�?EL���v+���F[l��߈ �5��]�Bg���;�\�O�^O0D�R~á>��+�\qjO�9b���D��ۈj4�N������.�a�'�'�!mx��5��o�!�#1̕u����d���~� )p��:#��<af�,t���4�7�p����*J��@#Dd`���L���h�<�;y������
mx�
-t����ᓻP�.��×J��ڝ�5�8��	�7�_[�/�����nrѧ��'�4�% �6�6���[55�s��㗄����C�Z��|�*7y�����|j'� 4���@���۠q���un���bd��o^^��~��	�9�Z��`���S66N�-���4Hb�3�^����i�ysV||��vF�D����S�Fk {�\������^��i0���w���y�5���:�l���т��j�vP?�|>�
1��RRV>+nr���,��4 �&/��%ke`p������i~1&%ZE�Z�#����ȸ��A������7Y�=:_�?��>k��A��
5N���&N��w)֟���Rڎ��k���y?�z��Eu�%��5���/�ɭ}[8M���m\�V��)�g�ٕ(N��6��PZ����kgo��ZM4��mSA�|:��������U�D������χ˜붯u[�p=T\�����2>&BP�O5��v�����hl8�Їϗ�����f9��de�HI"���[�����*�B�w�n��Rn�;���˷�~�AP�,ec��;wNP,A0V�.�s;�|��\�:UM=z ؐsެ��r0]Lv��W��9��=fp �o�1�ˍ\ɭ�~%4�b�E�CBE�p���:⏒�n{Vz��w�!|
��^��	�~�U^|D9�<��k�c�*\t��q��f�W��٬�UX���1�)=t�RK��e�go̓,���q���ӈfC6�(���Ysݑd����yӚG�>Ix�|'!��^�|�?Y!ގ�ll����	O�u�W>_��dv�D)�W��
;�$Hs�����1O�%�(��Q�n�f��7<�75k�U��Y}=��s�>�H�F�'Ҭ���b��������9�6�e���<��}�f5�����z��Ÿ��[H��Y���85x]��?`5Ŏ +v�S8�e��\B)��3'�(X�]ܢ�hϼ@mU\��K��Y��d����*V^�#-����~fu��<$��������6���oL�^��̡D�u[��݀Q���H�Zk��ڑqů��!�A�"�p٬���B$X������N�#=
"/�	�j��f8��z"V�)1�<�?�9P�
pЅ�G�̄>�1�����7��@WQ�hB7�_(<�&ݟ�۸���ͦ'�>�����]N�� �����v<t���3�I��/��bp���ڸ�zd����q�C{(-�^@��r��r��!v��#��}��o��v�b���/aF�]L BR�$��)��X@�p��������AG�@ੱ��ߨ�=
�qմ��-���}����_����4�l���%0=��-�	���>y7��ʿ@���=�8ΰ�j�dJF27iq#L�8氻ؘݳ[)q2��O�L	<���G�,�M?=��-�ky|��lM�H�H�3�	���%:cX�r�2N[A4�����>���S�y���'-Î�����t9gK�ǨI�
��~A�_�*��`�0�P.���E�T���2fg���X?�a�Px;U�Z�����>��^B	�E���|���l19ě������C�,�[�לAz(B���`+�9uZ;����f��S`����B*h޾Y�02iI
��\= \d(�9mV�)g� ��S�=���\>D"C7�H�U3#��q���$6D>fp��sTV ���4eV�?��"�ر$���ŉ�	I1@�H������e�}A��w������^`�,Oo�n����4)j��}��S��Mcc�q9i�y��a3�&&���V�N!]>d�m!C'����p}�f[�~F�O����?�e�}����`vd��H]"06�2/-Y~�
玾����hv"520�2(o�Q52�Z0sB���1�S�_��A�(#�/�w~��o���?��j�D�8He&�h˛.8������a��m����#�BHX��D�# A���>ǀ�{�������ȠUP�ua�]#0����S�D|���RlJ��s�az��)I�ߌջs۬�U��G�mt��/�w��2>�P�������'��T��I'H�����=��_����Z�o�Ǌ��k����A:)�	m(j�����ł߼2�uB`�}�瑅͆�L�Ѫ���R����3`!-d{�9�'��n�\V�4����EO<�T�Q��$H���� /(\%DĬ�Oa�`D�RY��T�(ʝ�j���&��WX ���Y�K�J.ê�i9���]�{@��B�Ӿ�� �(	�  ��4�p��x���+ß/nsU��"D��67��.1�j!0@u�Y�#�{rm �"S�!����� �a%���@���."�E��D�� Q{����'|��em��@�����	������e٠7�	�J�j��Y�ŷR\K�zQ]��X�}����"��A�S�nu�%�缐֭������R֦@�kيc㽩x�� Ah�lS���h�6��c���;��,Ȼ�	|�ע|ܤT!�/Q��1��y$e�!	fB[pM��}
,@��5� ���&��{�8��5��W$X�㗉�b|ܜ����+/�q�Y����3L�Fa�������Նed.�j1ό��p�|�Q�_��kZ`��O����zH��6/�+9���~��,5ۂ�<GCW(a\�����#�xz����6P"*5���b��λ��ȟ�_W���yqR$�T�Npi��[VV��w��N!cjxG�dXP�'�����<~&̚{����_�.PA�<���J����G_��7�eVo1�?L̰�g��,���oW%�<{�|����b�*޿w^1�l�������l�2�h�Z2��US����!:q��L�G3�pW�sz��u����A��Q����L���e��8��5%EQ^a\�}n�5��O_G#e�B�l��S�UH�9��>��y�@�:��Ϙ@?B�tHho�3��e0�ѮK� �Q��#��n��(�)T�4׼1�Q��5֘M,��o� ����I{��s�L`�{^z�#���%�Fc�� Ra�wo���(s���E��y<�!���	�늟�P��ҧR�c�ģ�W�O����~�AZ=.*~��w�ga��X�(F)/A���b�fY̛Y�Ӧ��pؘ������0�f�y�h��i5Jiz.j�R#���E)��a��7L��D�����Y鄲s)q�{#+��"
�c��a|��#@��+���e2��
�N��Y�ck��f�J%���
�L&vX?Pl������gr,=�f������ȣu`�l�z��V욹��О�#�oj控��Ox�2$Q7� �+ �] K7G ���.$������yKht�z��<>�U����\'�8������<�I�HP�`�1�<�X�
������xl��ag(�!�wH���ڦ�\X�����b�x��Y ��UD���F[Gj���c�k/ �ڒ@7�Lf�,1HX�kw��>F���i�7�W�k��@u
�g����o9ߑ%/wzR��M?%q�_J5o�j��_�ѐ_⥏�'�EZ��I� ��if-�t�s�E�B�l�������.�?����7�}qW�yy߿@`�;��U���{}8Rjp�X��z'eA�f����~�N�S!)$}}�O�+B:w~��wB���{����,�=[�V��:�T"�7�pYKC# @~��<����1�Œ�'�	C1�wA��ˠ��.*x�d��/��$w�@b��Ak�`�ȉV�$UET�ܳ�
b2 ��ac����>"�4��ro��D�Ħ=�{Cr��#��4�il�	�pl���F�1V1���*�=��?m=������=dز��e�	���^����:�\��N���������<�UI��)�HQ��^�����!�=��N;)��k��鵏���0PKzx$a]'��-!-ȵy�˺�-V������c��}�vL"�8���	�'���������6��v�O�6ҡ���o��K�I%�kf�n�w����L��f3��tL?�H�&#�~ ľ�S�2�6�J7m �i�Q��)�㝰Tϙ�eB�2�b���ů�)ύ�^wtX!+�jm3&<����fw���6-h,l.�͋�N7^(�����p���?��u=v�[�rV�U���D��n7�CO������d�7����t�qs��>�{� ,P�hc������%��q4�������"���X���T��O!l*��[;?��V|���.~��:�o�s��c.ĔY�I��~L����I��	`�R\�!ɍ<�t��!#��0Ւ����!MCC1&��v4��#
W�8ʓ1���0���c�}	<�X6���#6������բ ɂ�o�䢥�NO�S�ɫÑ2qf:�����ސ|�H$�'�c��g�S��ne�5������I�͸t��D��xh���Z��d��O���o(�A����Ź�ދ�����hv��N�%�jxR�7��(sHRM�����:����������O2DZ2�&���A[�JXHϹ�o���^ǚ�d��E��Y�c���炾�I,�� �?)���[�f�8�3�:B�+(`�U$`��RR�vYtf�E
c��.�J�n���Q�,�C���:D"��e�ViF�/Q��V���yFi�5��]8r1�|�9IM���A'���@��45|h�P(<�fϹw�OE��5��Otn���Ue��b���2�ho_��\���k&E'���W�Ĕ�~��efj!k*���馯�D�:<�p###�[|���|���k�E� U�&�(ʷG��pa�j&S�0�=<��k6DP�lZ
AEEG���O.@)�����)�<lrbAPrlă��o@� �2��}�"�M�{��Zd�-IG)�G*���w5A�'P����[�{��,�t�rR�E�?%W �"�����������}8v�B͙ 3=1�˗�Ђ��	G�%�`UbV�o�ҵ�BW��@��ۚ\�џ×iT�tf�B[fM+՘Zx�0E�glZ@<<T����.č4HO�K ��9X�@T\ �[Gh�%��FT�r��Y���E��g�s2᥽�%9�4ݣ��2�Bb���O��`/��'t���Ƚ�x�)�w�S=o��Ӿվ%�y0�U�0���pp�C�>�3C���_��T<y���#���h e�F
��3!z�� YY���hx0%��*z��{|Wd�T�!��kg���#��d)�Y�w�|�l���DY���;uOf��N4�uA!��I�d���g�ZK��ڰu�0Lc�S#D.�!��~>0��M2}I4|b�ɒf���9^A��d��ǈ�"{�`��T�[��E�^�L]&֋����S�?��I�")�P-ӵ�и�|�����222�3c�Yv�V�
2������R����1���X�a����bϰ�zB�~�FL`�'���K�Xm�Y��B���8��-�͛?�8m_#����3%=4�E��T�]�N��_���V�m��߼B��xv����{����{Ńa{��xNެrWT;6� �r�S�����U����>eCAtU~�ST(+Pߗ|�W��k&[��ů�3��\��#Ԇ�8zWQ\� R�����z�>@@Lҧ �+�{e�=q'��yB�#6�.�;��FG��fS�+��)#���wn�K�}�x2C :{��lZInY!2\�e��[�R*��� %��,$F�+9nV��c�p���<���9����Peљ��v{!�9��W�nd���6���O|����� Cܮ) 6�[vI�#L#��0`el�L@i��y�UڸЧ.��7�H��]�u�[�����-�l��L~ ��mT�$MQޝ���=�֙��Գv`�Q&s��a�M$^��}¤��e�q�k�=��%�p��/2��$Kp�
�$]��cU�8��G�[吽` ���BAI�'$�rLe�wnpL⧊,�>�Q����+�pGB9j M��K?ӄ�ή0B�s/~�1������s��[��!�BC�@�{�����R�*�w��)��B�t�"G{/���B�M�>/���Y�u��7���L�����K9�:���({(�|���Si�GeF+��K �bb<����X��ө� �#pSX�G�&?�5MJy2`���l+�< ܢ)��������Y�P�0c�U^j����	q��XC��J�ps�������=���s��@�숍����	Z�6�w��ت�����O$�#����ʔ�7����(�5 wܸ�b�!�b�q���D�
��L����N]:W�hA�phpx:E���6��J�uС��0�6�KpT��0�'Ć�1�����i�!�ϔ���>���RNp6uĕ�jj"�X	ǏW����#Ӎ��	�~���۠!�3�$��._&�8g��jK�o���2��'�"���ζ?+\�QJ���8jx�h��S��+4�d<��<lg-��WB^~�d�;*� VbǄ�)V:H}ZQ�b�~^��Gʌ3z��7�ܧ�r�bel{ftl7E�dDثpՂ|������ARj�S������ue��0��n6�[�H�K-3f�ƫ�O��.Hs��W�7��$�4Lk�tetkb�y`�"�/GF�L"�棂�u���A��+�nO�������a�HN�zݑDdQ��"��V)�?��h�Z�K�s�H�B��#)��W�g^�`��U����'+Zf�ᔓ�k��o�f+��Y)��0�p46q���Ϡ��z{/�6�֮r�Y������[�]
8���x�k�[Y��IrPt�-{�b���ǖ�#��κ4X'@
����ɮ�Ƞ�Pq��*t�2)�"�'�eļ�@t8]d���r�u [����쬉���^v���	��1�N���^P7f;*���j��Da;�=�=��0�G�A��+�g�i�$�'���#�[hj�-g�@�`:g�z����˜��U�Jy����\�nN�ѷ���U�����iJ�?e�*C�~��N��Q�P}�_�����@��V�SK<��]��S�Nh�����Z�I��z����P�HB�'��nw��|w������}��o1��ē����D8��b��W���dU�����~�LW��-;���T8�`�6(��LK�+����*����'L�:q�%�x���\����uS�M�!�m����v�P��a��Rh�X�8�殽!�C��ݎ���)ey1��	�����r��D���n�MFn�wsl�V.�<wՒ��Bw7�Dl�b9��i���`K7H���X���;��!���ȍ�P��6��"..O�H�v�MI���q�>�,? �Q������@���z:ޣ���O�����"ƾ+pJ����⧷(�a+�3+#��=���?��Z�M<���f2���x�|�UN-��߹�/���'r���%w�ً��:�^;u ��Q1�,l{0O��R�1�6��\Ծ[���{;�cބJ����)t"l!-�l�Io�pް�z�XrUL�*��4i�_�����=��5�q��Z2�)�1R���m^�j��D�p� �f�zr5�p���*�>����k'.��:�Mp�q���NA��h0��bļ��-Vݸ!^7k��_K^,� gU?�u��.(�b	�W&�:��ǻ������{"�U���}��3#�-�*�5Ի�����J]h���[�`������YWs�wW]],�Z��7���\����x{�qb���΢�!v7��r�lb����QnO(��˥(��dR�����!�?eZ�>y�6ddmr�rQ�*�t�J�ŭA�#��.YgF~�.;h�?���%�R���d.�L&��( �9��I?йQDO�}~P�z�#׮$�
�ȩw�:��+2ɚ��!m{�.��Ԋ���p�SBݍ�e�����sn�|�p:B�O�Ͻ \�
D:�|f��|�ee�C(�<&�2��{)��q��/����x��(���%Ѿ1�kX�ٳ��a]���p~vO�I�zT�݇��{U��u2��L^ �޼����kl��t$��N�M�%�?�+�"M5q�s6�8�������vB�$]��9�@SW�(��3N�^q�{��/_N��oX3���~��Ǭa.�786(�)㗗�ݎP���jH;b�;�����D'{`@@={��^(V�U?�q���sit��p���[����i���h���$��f僗��^m�T�a�G-+$\##vÎm���S�%�2��]�m��9&�����hp\DC8�Ћ�B ����>�=���<�����݃PJc��_�В��:����YKn����3�;_ҼI��?�_�N���v��HV/%M]m�6���OO��/�:�	0�*�k�z�Mű�{s�;,��$i�5Z�6+;�wi����:7�_h�E'����,���K`�9
]�
���.`=��v_�(���ls�_���ȴ}+�=PR�ʈUzjm��4��� �#ױ�Y���O��F��DJ�\�Me�#u�\��t����2�4u�	Y���(#�(�v���_���	_�$wb|����}��Ğ�����7c7m"�\l4r'��2��\�q��wysr2XC�Ws��DAJM^n_~�����x��<gy�%�7��pki���& ��K�'F;���Pv�ʰ�����h��Ù���	
�������;�oI�GtDW���@3�����)uwt��[@�ϩ�5^��L����}<���(7�T
�K%Y�d��r?�[�y&Hߢ���9t[(�
�%�ޙ7yF~�m"��=�yRi#����2򧥟���}L��t���Z,ȝ��~a�,�q@�=N}�����I˄�_6=V��b��t�=�{���0�;�a��佯]ع(>+/e��M_$b��N���*rm8��乪#^���q�愻�#�hO�9tX�l��m��I��p���F�a��f�ůL�o /Q'��������v�bV�Wa_�o�}�Ӷ�w�/N��$���g޵���a�����Z��M�XȘ!*1��ܐ�?~\�C�g'<\W/��aؙ ��vmIj��es�#�G��J45�Ii\��IQ��|9��d��I����:JyZ~�y���������7į��Y:�2O���o�[�9��6X����r�����X������"zlI6d����^q(��u� e�<���فrk�.Z�����p�y3qU�Fܦ;	w�O����>7��*�L�qM��p4�0�}I+?(@{��x�����z�(���$蟺o*%G��p/�㗼�al��/��=�����R������\����kA�0Y�B�zj/��o���G�ՌU��_P���7|�͵OU��B�s˞�q�vZ��M���R1He��tw؞�WI�S<�K��~eXÓc�H۳�?�C̤J3��a-�B }�N�#�uHx�$�9s��8�;�����[��K9�Stf�]���_T��t��,��eee��o�m[a8�-��I"!�w�>/���'s�i˗�I��E���e1̠?٘�i�r��XS����6\*�	�Q|��9Diu�W������~��fH��[a&�³��Ze�s{	�����G9�����iG{�q���J�p�v<���P�rW,���}:)cU�R���x�b_r��'�I}����6�bJ[OG��Ϋ�ޞ�J^����U���<�"� ��H_�]�<)�v۫��"�e �A��1KО����\�Ia��;�ܡ`�ڏ���P�����'
+�7鮗y-e��#zz\��Sm��Ġ�DUkQ��g��
�g��ٮ8��궆"�.eNO�D�T�;Y���,���C�TǪw�oGn;!ٕ�#'�Flg��8�Vji�%B5�#�9�4���t+��{�,V�u�{]��M#ps���ɳ;t{�r�!�g��V��IȌ@�)ʋ��Bd��qz��o��'ѐ��0b�{�� ���4ґ ;�ٻ u��9i�����K��m��O���H�z2R'^�Ywr��=�j������Z� ��#`�t�Z��ҝj���d�3 I�. B�ַ:�/̕�g����Cwx�xJg§����t2�Ԝ�"\`޽<�4�#>�v\�4�d���E|Bk`����ߴ�s�<טIo3���ಐ�(��kF�0��������ny�N~���B�t��,ݩkA������VW��!1��M[�muP�U@r�Z�����>m|��i�5�Y0�k�C��}
��|론��|9��Ӧ%�;3<,���h��`����Փ�S'w��������Y�yA����0�PUᚐ��2�i��U���Ѐ���_�
 8mN^��K�5
�,�����ۡ(���6�n���X+��0OR�pl�M�IZ���U'k#|	_:����U���-O	g��)���q���x=F�{HDu�b�O�����d#�.����,��Q��,4�
�Q'J�4���kɞ~�X�b�\��_���n-��
E'l1��[�w�OM�¹M��,��ܟJ�s�Gť�*�~�?��Ϣڪ1˼p��|�����`l/��9ރ^�� v͔:@w����n+�)�,\��q%���hW�e�m.���݌��1�wOW�.�eg�(��
�]}��b������NLH������E^N�x��7C1�"��Z�\\n�RL zw�8�;[y�!�p����"���S��x�V�7�ca�� +�I��W3��\M�>���^!�E�ȣ�gy�`��>�tE3�Q��@1���l�C
�gq���͒��Nf`���^j3��/�C8J��Ռ�g��.e ���`?�y
Y��_I{���d��Ί���<a_��؝0h�-�Q>`��)��Ӈ�3�d/C��*�^ԍ.�U5W�5z�K��</�W��!�ڮ���L1h��_0��9!��GdM�U�k�n��d@���ǿ>��pQ�C�)/�f(��M<[3��h�2�][��?�V�˷'ޯe��U@���I�Ī���������)� �zo�&M�G���_}LMD8��߷� ��v;O�������_z,�&�� �₊*���:�c��e �q�He�El��3*כ��3na��k��%��GRvH�l�����5����ci� �� ͚�\ �0w�uƧ}���D�繁�rd�x���o�uf�1���ܽ�J���Ȧx��B�1zx^R��t�"fne�H�Ӧ�`Kމ޽�m7���0_����j<�R����|Ȧ�����|���7��]���T{ݏ��qB{cB'�����$�>�n�c7�@�[�8�b�}t�� f�;�K�{��)��ս�Le�n�p,���k/�������x<�+�`h�@h�W��Q-</���@�׃�.��ܖ�ڪ���'�8�d�(ｖM��칛��_i� �9��0Cӽhip�k|��4����`��ޠ얫J����ѐ���b�Ɍ��G�W��Cr���=�t@��5~�w��d�c�ZWW77�����t��-���N#���W�l����h4ٳ7㺥#����E���r�#]L74̴��e15��jqIT���zW�̗,�<}��@�@��{�F�v]]��p�p�Þi���	U{�>5:jF��Bd����L7�]yש8�x~��f��P&v_E=�e��wp$�i�}��ȳ����#�/g�E�r�YJݍ�����ț�&n������}_����H0�h�z�ۂQ��x��c��4��m�BcѢL�����D�U>zMs
�z���
 � �p�RĮ����y��~{��k׫��tqR��x'����y1��wC��'���[~��$���g�����&��B�?�[�TOO ҾV�Z.:���n�����L�SV�淹DA��6]!�x���3�����5%�P�,���z��]�2U�����T�?�i����;���F2���+]Senq�~�����2S�a��̃�n�Y���.��2�.̤�g�������n{]���f��P��*�ǎ�eo�F���Y��A���c�@At����j})�z�m�D-ۡt_�	�x_'�ϳ�$����n���S� ��
yyj.p��ZXVQs6_�o��h�d������z$�G���9PL�@��]Ƴ"r~��d��w'QCv�|����G' (������j.X��?ҾY 	���{�.�h�~��أ/�f��=F�+��Yxy7o���{�A���Xo�� �;�y����MmM�h�#x^<ǣ�
X(ґ*�r,��t�(MB�%x��@��B�RC ��.��"��� j��~���Aa�5�f��yf�w�����/��ɭ���um�2��y��W�Oݫ�˴����Ta�6��I;���Vg�L~AY߇�c���U�3����fՌ���� K�Y@�kgR����Ǭ&H��/��xd�4]�_�_�����>��jnƯ�3:K�6<�F��i^�cYJF�D��Y�����)֡�����K,GC�Q�=L���%9`�f��|�Vi�}�㪱�ε
��kLW�JW7��bj�fK|�u����m>����O�<8Yw��@����^Kq��zgk�lׇV�Ƥ�����ϟ��Oʈ1=ѽ�~�s�k�qB8��6���
(b�f,d2��s�<)�N�eLMYc?��Ĉ��	����s�\�KvO�'�ħB��[^��SY����ʰ��'����xő� ��՚���e ���<�@Pk1E)SBcf�6W{b�>tn}���ʦ��ut�Ts������:P�y*3��E$��td��t=}��:R)qv���8͠�/Ap���#T���
����8?�>���[`z��W�\�Ҹ٤��I/�U<B����x��$-~�
��ީF� .t�J�9	I���W���$$FP)���nkq5�����/D��t=�e���ZXo�H�^xn nČ�+y9���3z��lE�ԥ�͛
[�Sl��2�ޅk��j�W:���SiR�]�e�~^����}� Y����>kT���zcӹ=S[�0�
z*SY��:��U���BC~D2�ڒ���߻I�ۣ+�>2P�|�-f����$V�����U�f]�+�~-('���Y8�hO�l��ڢ�O[����C6��G�a�D����x|��؛��M@;ۑY�
��!o�Pp'�P���i���"$B��[��]�����bV��ab����iUي	�9�*�<Z��O�Gj�qJ��h%5gS��O�<�������U�͒��ǘK]>B��/���f�jQ�3�A��Rl��b��I��E�=[�в�o�R��/ަg��v"�r��U�$W�ߠ��>T)VQ'{W�q< ��L���9�=]k�M�VDn�O
M�-D.�C�(����AT���5|]�Jj��fH�4<�_]�if��w���*�8�_D��ux}E.e�B��ɭ���z�㜠ᠢ�;����b���q
�X��@$��Lz}ε��J�㚯�����n�F����M%^�;�N@L�Z�Z�Rں#ս���\��*C��P��7�Sg/#ϣ)$N����\;K���T2�X,�!�$�#�%�|�|��,Ĕ���&˕:� h?�Ӹ��Y�������Z�?�����O�{u/��6�#%����>��#�>�����B�)�'!��zq
u�C�w2�4���s�7�#?ǟ6�5�������9v�!�
?�&�Z���꧕O�=��I���a�yE��HC�'��k�dq����th���\d�v��j� Z�rw��k�(Q�������2��}�V��n��旮���f�?*����O�����'oj������;�@i��䞝�n%x��"&�g8n�w�k�7=��+}�/�l�|&3��O�����8��i�L؀b�[Lj������bY)��,]��l4�c�qU�F�C�Lv���D"�����������A3�g�+綗����ۙ�L$a���-����QOKJ�R�ɏ����_|L\pc����S%���"Ԃ��\.;б��:{���޲�g�\�����H��`��IΖc�:�RX��fPc��5V��I1��^�g��n͇44�b��������lfIy+@��B��f�p>	O2�g3��'��
!�@�~����-���?�lT@	�)猈�����l��r��"^B#��nMo�84U,
*_y��sH��Q���ŠzQ��}}�E��e��)�1��ǎ�PEܶ�!���S�WNP$B���\�������-���H�����F|	����V9Ϥb����GgLܟ4�y�w�����>8
1���mDR��kBf밣:�Y*�N"N�����j!�䏑�����+C �a�sfh���s�6L0K/m26�~"����"k�}���n��M&���ҙwex�h��Q�BC�ӿ4���:]'Q��]e^�TN�q�h�`���,�4�5�tS��
Ώ�{uxHDD$��/;e�R�]B���9�nfij���sZQX5�x�>a����޾��47"[�T(+�|j �cIo}c<����^P�$��riޝ��B�1�M�|mrb@��V��T B�n��W����M�g_(%�V�1�־\����Rqfw�כo^Γ�������a�����k�D�@�&�:�l�"Kcp^z馒1i�U$�$���@sp\����U9Rz� i^�R��WG�O,?s��Nuos�K�����3�<��49�~6�A�F�rS0�:e�c޷7c�Ѡ��i�|bǯ�%��?rF
\������0_A��:
.깲�N��<n��!Rn������2�E�*G*����
޽���ך}��V*�Nٌ��^l�����G^��L��H�*q�q�d��'���C�b��L���&�f@�E@������SC3�Kol��2{��fi��H_ő�K4!W��z`u���q]i7H�����z�vcS��|!�c��0ϣ]��g���)�Y�(������U�f��g+h��ڴg#4��]r��^9@/�^t�ِ������2�
h��#������"�$��\�����7�!�V����M��ju�a�ɷ|xV��E��ɩ� ll�f�Z��!��@9 !�\���v���$r�Hs���'�X��Q�?���_���������%��3��J�e�0<������KʫO�i:�%[��<�&A-Y��@z�f���+g>�?c���r�\�d���BA����L�����x�I�Ec.�(��fQw�;��b����Wř���6k  =��D��Ń����8���s�n��b͡?l�}W~%�ר3�_��h�H0�S��U���c�,η&�����/\�-���5��!��`r�ɋ8	�BA4����W�X���4�~�7�Ѳ�?')-��'cӋ�Q�����t1E�,j��V �.��~
Qt������� �afj��_�rc���z�q��6��9�	�@y�'��B�ie9���|n�� ���}(��sm�YN�ҥǽ�+���L��o����9d%~&	x���Ͷ ��R�vV���͍�;�M��8r��|�1(;���"�?Rw���PP:f�eP�@�^~&y�aS�����쇇��J��,)N�W>%��\���%^��g�Yd�����%�J�vz�d�S���`�,�i�I8M�'%�������Ner���T�̤]Mẅ���yy_b Y�k������E�j�l@H-(q5�S���UE>ԉ$�S��x_Axy��i^�h�*{���4pw�7)Z����{v0��D+�g7��_ ��4�o���M4�f�|������[Iq�B3�\��J�R��D-�,9����=mJ������{Rn����N�{��E���p�&4O��>mꁒ=�Pd���; ��tR	�Uט8^$��,s�8C.7)���r��I���6��\1��q�oD�F�o��Sz��(r��,r��Iv����f�h��B�*�]~*��+���=_�%H�R>OɜVl~�F��	En�G�"m��y+��'_�Go	�Xz=��jES��hS��%�\@�Oи�{��H�L��R����,1akѾZ�{"�w_�|�샮{�|���__�ʝrU��������|�����4���c���J2c�w2'zz�^x帇�1�$e�'�S���K����-�=��d���d��8���&˅��F�#����)9��\J_�������'��G��4�{�L�!K/v���7�_�7h�/�ɚԥ+���x�0�Pb�u�[&��e��ɫ�S"';S'��g�of�a��A�Oz�Ir)��z�|��{�������o���k�(!��u��m/b���T�d$���n >�=�c2YC��W��ww_���#�r-�2A><c���h_�,VZ�U��Ik/��K0�,+�!\�wҝ`[�0�G�
w�"�����[�8����U��k���,���&)%7@g��vx��==��ظ�S�ԐH�Sﶎ��E�A:�l$zLVO3��w��'�s	{\�e#�zN��\��S��� =B����>��f�v��_}�d}�xSxEZN����[/S�Q�x
���M����l\�����G'l_�����"bZ#�(p��U\Y����g�T�"@�=����W{#�,-�ў$/M?;p���d��t�5aGI�l����'�S+��[�=�v��
���Q�Y�8��	���2_��}��i�y�
���Ʌ>�B�xY����cB���f�);�oOF�}/�2��6r�^.���Bb�i��w�1CÇ\އ��$��sg��RvPZZ��2��h��1:ȭ�LLj�N����c���B0�:��s���]&��0���/9aT%�4bs~�o�����P�!��u{�tW��,b�}02D�{%��ow��ښu�^N���uͿ] ����.@�����4%��e�<���[L���5�XP�.����R�f��E��}Oa�~�) ��W��Oϫu)�=Pb�dN���}__йCh
S�����*�S�A��N9���N�Pv��H�3�(qX(�8p�0p0Imμ[�I�hQ�xؿae,+�����;R����s3��y�x���D�w�s�+?����n�Q��w+�_�䱢��$n��1rC�T��\~��pb��*��T���0�T#@"���F�sP@4vm�09�q̝�<)�qs�'��%0���~��&�/�����*����L��@�;����6X���}��#@�sP�z7=��RC��O�	I����"��3p��d���Z�	V�iFw�e�z�)S"��Rg�y"�鹖U�|
"Z��GCtm�Y{�!���|�t5i$��WE�%��:=�*&QH	���I��x����`��{�-ؾ�B��v1���k�R#pg�]��Պ�0��I�
�������yʂZ���*.k�=)���΅'���4y2����~�]���T^Y?��'����w�2�7�;C��i�>']ט��&�ՁX���P��&E�M�S\b�L��מ�Y=�y!#����eZ٥m'!�?:�����#�Π"����������}e:aJ�h`��).�����|풰%���Zo0�������@�U�8��pI5��Ͼ�T�gWj�m#מ5����]	�U�q�l��@�)��;��g��KKx�F�Vl��|r�ڭXa�? Ma����t��������g<�j����H)��k�u�l|B�����Po��k��f$s�+N*~X��q�;����!�q�S��-�U
��Q��'��O��
Y�C���%69*pM�X�$̫ޔ�/�,:�rzI>���QS
:�\�����:$+&&����Z&�⊔���ϫ��o���
/�������]�Y|�� K�́��������Q�� ��k��:�a��:�>)��wǨ�?�P���;�=[���}�n�S�d�+'��|�"
���h�7�n�w'�4�;_���I�R�k	�\70ܸ�\��3`W����=
�o``��+Qp3�����ّ?���|q��[<�Ŷ���88�>�t
	���IR�l-���5\Y���ɥ���.�݃ B><����c�ʫdը��+R�4F��-���]Ս�F�+��g��]�wW��/�9���7s^���]��t�t��������2�\�>��e"�Ŏa��B���2S���ȹ��M ���C�ڙ�8��07('��a��/26;�S�����?����D�.�F��wI�.Tt;�?���Ӂ��ZQ��A��n�`����=�p�ѥ�4ԗCB�D�iS���o	��+��S�����d��-��Y6�Y�Y�o��U`)s�d�����ۢ��I��!�K��;I?���#��N��Aw���V��h��"�At{XԕM+��4W(7������剋6�}�ވa�=Z=l'�v}�D���o��R������Uy�.(������ҤW�ȥ!NEL��
@��>�6ɭ0y<��0�w����T8` ��N��H�eOh����ǅ���N@k}5[uo�j׊���X�S�O��0��5U~@�"ԩee���x���4?��i���s1��I?���**ĴN8O�=L��� TQ�[ g�� ��2fR٩/Q/.��;�ؓ`��@�=�i��&U�T��ѯ
f]���)4W�'��ϧ�!��^BW��m�#r���)������V����)��%�s��U���[6�Q0��|�~
`�W�'Ń,� �r����Jw7�|�l8�yA.4b��J&��ط��(��	����ppH�X�2�W�~�du ;(�k
Q�B�~����)��sLU|��d !�P�W�#�SJ�S�@�p;�~c9�	jv��G`f�ڵ�kW���
jSԷu
n"����:��T���q�e�'�v�{��X�?�=��r�	�o�Wl ���YIW�Ĳ�&��,V=�+\e�9 ���*͟{��	'��!����LW��l!�M��*m���P?���,#;D�F�2T����L'�yӒ��ˊ��c9�U)�n��g�K�ZΉ�{�k9b^����d�s�2��s�ܷ�8����P���1���F���)9h���y�r�)RU�$���h�tj�R��^�Y��v�MG�O�J3��w8ry��*,�Z���&��7�z�_�؉�| ��@�%il%����u�M(��8<�('�,��,�-�v��~�h9g~Y3�+0���JX;]V�o��s�c7���`�CZ�r���h�UY@#Υ�)ʆ���=o�nrO�ts��s;�Y�lN�dS����ɸ:g$�8���י�nk�؍�H�.�8R4��G�W��٘G��ߋ�H�%�VK�,F�UA]�1��R�����.�����l�ƕק����)�����W.G�s.�Y�w�L�8;�s2�t�=G��d���﷧/G7��z�rD����
��k�|��6��Vu�>l��#:�r�X�hȉzH���~�k+����V��������ߟ4Y�ٔbqy�L���;��f�*���S��i�� z���BW���w��MM���\���9U�۔�kb��,#�18<D��n習/����ç=p�:�2iQ�k����#�Β�=�����4�t�u���
�P�Q�@0C��?M���m���uw���$uŨb�V�ۊ_(r��P� 5Z��*���_g�:^y��[�Mw�Lэ���TUe?�PB�v;��jCs�9�z�]����h3�CW�@��M5���������JT��\���
Vo��X���R�~[h�`�Q�����l1x�@��[�m�4���	��������2z��Elm�(�$.��s��"T�/� :`��g�}�8���"ˈYxRSӡIx��r/	K�)x9�ڣ���-3�}YWegËP-�ve�fa�n�J�T�rC�����)��U/�6ҕ��aS}$�NMN�GS�؜[�2��\b=':�z���/��gchUE�U53�|�x�RO^Rd����Ыu����Hܝzq#B���;U�(��h�|�oD������逩�de:�N7'ڛ��Z\��Xq�(�����~�0]�Ê��_��2�{/�'�|2iH�i]7���D�Ay�����ϗc��r	�XЯ���{%�s��{*�֏�v��=��uV:��;���;��:Ċ��ˑ�c�EW��N[��y����MJ�Ϳ��e&�^~}	%�v~���e��S
��@��@"�3e*a���>��f�D��	�\M׽�'u�"����,|ۋ�1^��OW�Si�f�^5G Eǀ���/t���G�$Zz�������2,��[B�����3��^bsm6|�l�����v� ��a�|�Q��%�o936�N%�<��me���4LP��v�L�=ss��r��(����T'���|�}-��ԝT3>M7�X�*��B�ŪJg}����f?�>rV���K~�O��^N�S�5q�U�>[xOw�O@������m��>x�����8%9��o���y�d�b*�$^�k�����q�u���Y=n����r�h=W��@^r��l,7<Meκ�漑�,-vGk�4��o�n�������	\j�&&�S�'��[9�d=�$,�q [ʟ'&�[�k��B�_�kڮ�J�c�-a>o,�:�w�u��~O�wJK����~*v������Ԋ�_b
�1iI�|�$�vb�Z@�VS���>��
��u-�HⱩϕ�G)�����g{X(xoLn56�����S�c_����Ba��k�f7�N���I��=!�Z�T���#����R�g�M9�ι�5`<���hdqik�5r���y�E���h"%-u�`����i�_��*��4���j6��z+F����EW�u��2?�̅U�(�uq�*�6��`j�z�=���򞈿��K�ʋn+h�A� ��c S숖���tE���m��ZcA���ٜ��Q��!��Ό��͟%w�;��h��Gi'v��̏��$���d2*�FZ���	��d��e_��U�c�L�������Z!3n�e�k1)��E��]/�����)%�֞�3RQ3�S�$��x�{C\���F���4됁�¯���:s<�e�����ˊ�A K�Lڳ��J�ۋ�Qa������ЇV\n��[e���D���J���
�!w^�^�Y�Ў~։�-�PJ%d�wL�n?_��+�S�r��1��%F\p��?
wEˠ���@�YA\�x?�V��2��sF�.�#��0��E����W'\,�>�����_w����8����[-Ut�e��]X�&>N�-��Z��#%�*��QJe��)h-=fQ�Gdە�D:e8�������p�H'�X�{Mo�3�2�\�-�|�#��Sdw�5��cG����M�X�,s�Ƹ�^���B��rRU'IDK�VL����S�Ů�ʑ�4���_��zA�5����,p.���K��+ʅ��⥟���+��I�$��:z�($�z_S�]�\�oPl������أ�%��-m��|/I-���ˎy��uJ>��Q���i��]>����IC4�l�ԝ����L��)�7�]HY!Ng�6�H=v�>�1�S��J�F�T�OV�!.�p�hc٬r�1�c���E��D�@�Bb1��	���;�U�-//|ɐ=�y�0�����=�[����Dm2�/J顔�TNw֫6��y�.M��}��J��ܺ��7}���9��X\Q͵��������8�#�ڰ8��:i�F߯��^�NFU�f�X1�%J�}�w3:�u���\����!���V�����h��O!�T�ĵ�x�dsk%��f��f�t��4����dDt�Vj���BpיrLkk-��c�"cϽ����ٓ�B^���,C�8[ׄgk��Z�FsT�j�l���!z�E:0[.�4W��+-XxB�B��I���&�@��%���6jZ�	;��e
34A�M��{[�X�;wշKG�/8���Ҋ�_f��0�a��X���/޼�e>2s)<���J]�]��?>��&(,r`��)���\���23���פ�eհ��6N�}�*d�����	�����=J�;٢�͆2�"���m��"�""n�̽㒶�&��T��$S#�I��8H��1w�!���!c������1�[��q� ��Y�	�s.$I��{{��VmKv���;j❓[��I�0���L���r��e���?�<k'2c�sW�����x�����J�xa��^�l������%ΛbJ��f��v�綿1�d?�A�R}�0�F�k�~�pW�)��"{X�بCs���y�>��๾�t��k�3�ƽ.[D��y�Q~�LGr�TR�K����4�}�%s��~�}j*��+�1Bg�rf�
-���c�'�������=�������E�Z�Ԗ�m[�SӼ�"�VrR1^�Q�n����!C��}b`����Fs�Ub�f�n{��-���XՓǎ�N��v0����Z����f2ʻ�sX��*B�|���ư����H�;�dkTs�K�'�j�5��uj�`��?��˺��C�%�1�]3���A:�ݚ�~��#���N���eY��]X�j�@�����3�����)��:�Y����	��7�T�<O���"�k��C[��\_�f53�.�eco��z���n��9Z��>�925�X��5.;���Ǡ�ޫ"��3�T��K��e�n�b�~���wWR&B�&2��Ѣ�S����7[���_�փ?�����y{(�G�)p��`K���bk�Rq���X�V��>��э�ޟ�P�߬�Y*��h&�	�̿i��9@����^
�Ԍ��KYN%���q�p��4�mw�X�\��޻.��9P���+إ\$�(�%
���m���҈7eb�qxԦ�����^.(b7�@���Hܞ��1�9H�i�IRz�0꒰�y�t�����Rz:���v(1�����m5N����L�_m�0J�b�]��Vf��Ւ@|ޒ��%*+[�i��}�a��B�3yl�5�j�����'��W�.�x>�]�l,��M�t�er���"�5'�htKQ'�r�d��N3(n�����f��+�a�ξ}l�붟�g����������8\����魙^.E[Z�
ڡ�|��5}�cl,U�u����E^E�s��R@�'��F13����e�b$�iM=[ٯe���添�ˌ���(S$�$�)o��f".��>@H�?��uf1�T [���b�?]����ѨJ��]����{���2!���5�i2�>aR!&C��b���߳9��Hqi7N^4��.y���h����c
�|�!�?z��1IkiIYm�|�[��������HlM2ٳ��4�� ���+�-�c��r\��X�f[3L��p�;(bv�kavQjT���ǻa��!���a+����[x��;��b֔�_����՗̱�x��v<��v���\D�j���xg8�d�ѫǚ䪃�q�����>���=Yb>��B��dX,��[*������A��v�莨w]��p��ǖ"5���a/���[�}�Y/�3��8�FpfN_�x�;����&�_K��d���᜚��	[��E?�=����/��6WN����UX~{��rw=v�1Ps����h0��i���d2*�u;֮����B�vߏ@���K~�U�i�U�Io���%	�'�D.����A>8�p�	Er�%>�~4%a�YX����G�~��mwд���i0K��Ihzx[xRќ{4���OV���WBn�X�z���,���U2�&��2�ɸ,����ڋ�慅��ig���f�(?��*v�y_4��b�n���?VF>}�rާ<��UH��Ug��w��R�"T�'qT1C�jI�Ӣ7�ʽ��ߖXqkQq��D0:X*��봳�ވw�����v���Wq�WAnr��aC�J�g&p9�JPF����Ut�+�������F]�SI��Y���&��>��7�m�w��M�;�%�R�'��;L+쭧�$Ó�/�mkmM}����'��^J��\��d�_Y�V)ݕ�S噾�Ǭ��O��A��;*��C��c�~|�	j/�EA�֓
=n�c<<R��rH�����e�ЮP��g0C��n�V�o�������-*������`�l���h������B���8 �Ǔ
7�P�5�Ɲ�������=����Vf)��4�������~��G�~ :	��S�ʅ��XGi��Y��h�<oꇸ�=q5��1���F�GF�����������C,���.]��'�Gc'(m:*󗹾�=s����ܸ��j��wN��S������Ű��X��/I��	�0�����r;�_Ɍ�&d�8;�~y'�)��ocE��;���?=�rvo���H�t;z�)s���c�D4��J�/��@��}VQ��B�ʱ���7��E=z3��ٚ��8�H���a.�޶fc�5�E�9���%��8(rkV�s�X���cJ��Z��~zO���3=+ l�ԝ��c< [����j��辕LO��8�,X����r�B�u�u�R\�fO�z�����sf���B��{X�	��!��G�U���E���U��f��mDf��5�Lܽ��/��-5T��o`�t9�/j~�h���-
��΅��z�pv,��4V\�����ffl�4��a�Y#��1��s쮀�C"���s�
Ųm�M�Y��Б��9]i��"x7|�r����w�]���������Ǽ�������������_O��U��-�=G���E������N?$�ȯ�3ʧ���bk��}�i�0"s��o�gu�obe�CoGE�4PI�A�t^��vo���wv�hW�a�!�?�5�CZ�Mȍ�[9y�ćp���lTK�v�$1�n7���4�*�Hqơ��b���J��S��z���)wo����&&o>�V��mf�f�#G50�+�	�q��G񲃚[�0�7�g�M$�iD�<1~���I1�w����bb�d�E{*��*E����Kdajxӱ$N�p�,T��őJ�J��g|��:��rx�Z�ƪ���*?�հ��l��Y��;��ZFH�D������n��[���͟.k_�j��J_��#\����G�/~��9��ymӚ�7`�6TV7��2�4����N1{�5��JL��#on��kj����ᡢ�&�P��*A��³Ғ�_F�|����\�4R� �;��@"U��N?�I��*�r�?Z]ɸs�@�����>�F��vt���Ei*9�TS'�0Ƌ'I�m~L98$7�TC�;��{�k���r	M�Wlo���pH�j}L����l��	���c����|BT��b\)��װ��{V� ѕ���^k�=��_�AQVP½>�RF
��qݖ-��ƨN��M�]�vJ�"xX���P����s����ȁ�#�/fd�p��P;�S�5��	���L�[�@&я�,�t��D���0��mDt��!�6�W+������S���^��۾��\�K���B�e9rP�7���$�*uh�1��GC��]XW����U�Y����@��O�rnU����r���+��:X�e�SJLWcc\�I�S�8zǩ�f��W�B���U|[|P�q��90rV�x-*��U��n�J���/ݣ�}��:�*�ۉ)_"j�2��Q%��+��p_#Y�����R���+��	��hu7�	s��l��a��(a���[�K�q͙z'��>�c\�E�<^�1I�m@5,�18U���W�-"hϳ�r7m��9��`TI&�p_¼�����<e.���:e��
"ˠ�jF�<�4M������F����B��/Csl0T)Y�_�]ϙ���h���|�d�a.������;0��_蠴��8���L�\����:{n�L����]Y��.W�Q�k8��&�A��㼴�[F��-���lܮ�����g#���CO�:m�����e}��0�|�jDf2'h,�w݋\)wV�:��mo�b��~�.�[<�m��5��$�0�-�@�>��WH�i��.�WP�8�b���l������f����1^fb_�7��5=�A3D� �C�����#��K_��ǟ����ۻ�\<%3C>9bCo�mˈUI%̞E�_�Wu�X�G�"���To��O��VP�a�A�*b�"4প��-��{����D�r�Q��f�f�!���r�DH�j)P���_�E���T��4�9�̩����!|+��}��L���K��>7��gI�O� Ύc���>�q I�kػ�s����\w�w�}�EUTn�r��S����$��m���[�T�v����Sr��=�`���MO�%�oU��̔0��y�2E���[Y)��JU�o'���:���o�4}e 9����X	)Z5|`��w�^*��M���������0R91����;�{��_����
����t�,jt_��Y��A�0�a�B��r��+���L��l�1:Dm����12n�rg� �A�ۿ���|ퟩø�	>�$�M4I���XDp{��:::���/��@��{c��e�U�K�c�ۛίzk�v����9~�*�&���u�F�-$T�@t4�F�cd�BoGO^<tx%U�VI������3�%��2XX��Rnm�^��JM��Q��jȃR?u
f�)�K�KuB��#�����݄O�/++�}w�[�ρ�A�Ɖ��8�ǰ���Q�0��V����)E~��E�з����;��Z�0�M�`$�"�x�e�tu� �V���a�h�ذh��s���W���N%�о��*��p�c���G�H����Z ��"���'��}K�0�(%a�Z��uy@������
6�H��\_���?Tgdd��a���C8���p&�+�MX�[�׶��}��\���p	��[����= �=�!�,%�
4�ˣ8d^�5��ϛ�,���V���"��1�r��u��-F�R��{��Z܉X��*�Ճ����}�;�po���\I��g�)���������RUF��"��Bㆱ�è2��=�_C����Hs��,(BNz��Ek�4��ٲ�h�‐�J���.�y�꠼v���F>!���#����V��L��ԍXg���!숗�.��$��Hռ��H�	n�Xd�9�r���m�gЧΆY����;}Ō����-(D&��:�	U<Vg~��n���{χ�,v1�+�5��*�(,�0�/c� �!ܪa�5�Wb�{��,���%���.�{~���-i�ְ����m��xZ׽,��������_�V�[J�Q��rN%U����Z�)\o��R���ZC�>�9Y�����Ǉ��Mվ_���WK��ZQ'M�d�}?o0�?0��������ʻb��s����	XZ'ki."����Bw�tu��5��v7�H06�c2�4i7�q������3��m� �.<��<�;Й�����C�ɁZ�#FK�lP2Jv��Z?B��] ��k�(7�ɡbd�Bm��:k�Th$��8�L�)N�k�� �Ĳo��[������7_�&�qI`�g��ώ������j�F�'�K�4��Ƞǩe��22Pz�����|�O�RQ�G^�tčZpuD�$�̾�on�PL��2GG;8׶H�JGY@ ��4���4�;Mu\`�V�$:/�Ý4�f�J�=������Lk��d�5�uվ-�p��%�LN$5�E�U��bϯ�ӛزՆ�gӔ�J��;�ƶ�L#���m�j��!��o�$�_�Y����b?PT���8h`u�o�`�_bYJB�i�?�9.�\{�tw%�Zx^T��;7�(j�{�
S�Fo;$e'�$���I�QOi�q��]i/Lmmj��RgZ������k�b|7���KLz�m���)�.�ڂ�w俿H6�K�y���x@ZC
��A��,Z������^#c�;J���*|:>,j��	�3�Q��EUMr�0/�}�9�z�ϳ�$>>���Ϸ<El�0��*�x `Ƹ���l�UY��@�c��*��岾��3�-����(Ki��1A��z����G=oG�T�2�Cs��g�P �<xS���|N<�
!L]��oV��V��<��)ϨO��a���m�]�� r�'�F?��!�8���~FHXQ=} �s��]d�,�c
ך>�I�i��990Q�V��t���[�.XwSV�$[^��8g5Gdn�*��_6��)�Sx��B!���L)���S6q������"�>�v�vc��)����
z�����f}��&O(�@���J^��4����d����vҏ�u����k*b)�u��elD����ăhO��㙚�b�����̕����:�Z�(��R�&����g�Է��T-�P�9���F�[��qf�	��ᰂ�p�
�ж��$�;A���ˇ�=�U;ǗMc����uהX�\*5���I;#J�2�z(�i#IQb�]C5lQ���k>�k�g��(iFҹC����
��pN�7Y���Em���70xM)�; L�^HM[t2�1M�K +Q�C����Z�E4^(��̦��1s�?-&��	2/��F2�M�<0�A���&	������wu�y磌�R�!��q}-�IC2O�'���tW�z�Q/neU"����p��2�T=���Vŭdwk9��>@��(I{?X6�5��OF�kD?21[���� ,���RRx
u�2]���Y�y�$�v����XI���*��|\³^�V��Aӏ-�e�IjJ�o�ȿ�)���5lv_�ax�VV
�Jߊ��$�$1@"�p�{OѸo��T��4�O�^\uHT�5�T�{��<-~��X����vkP@\�e�:�ފ�v�b��o ߺ�>2�ٌj2��d��ET��Q��'�$�������px�(�(&I���M0�ǅw��Z}��kJw�p�m6@��X�+��J���8&�X��:�%e�0u�{�Vk!�`ySоt���]�9�=��+_�u���"Ҡ
�0�ˉ�[�sK,6n�	7�8�a֗���~�i�1��Nw�~�}����Gף�Չaz���ݢ��O�Sfޅ�L��B��2%J�c*�(U)u|�N��_�m�1>pb-s�@�Iuz�4���~sm߶��afs���\#���Rm�w��M<J�K��/s��qB8�E!r2��,�a��}ȑ��1� �*!?v�ܙr��	p5�))�c��$�|���'U�V��Ҵp��Ju�tYOO���K$�u
��c���Wf��*����'�I).
�`jW�APS`L�%�dXK��[�U�b#^�P�}���M���t�{��1화��As�F.�ݓ ��������|K�kb�#��m���=���K����]�c�_�mX�^��0%mz ��L���r���x.w�J<�c݅�b���22Z��?��19�YQ�[��f$�`��I�����!��}&���]�Y-�:a�beͯ�����|Qnfj||��b��x�f��h��Ԥ98��Ql��zmzg>������#�ǅʱ�â2�eg���چ��|ô|���2������m/U�s>�޺��a8�t����^/��vwc��������GyOi<~��D��k�Y��n�.��j�؋�5[|/��zL�.3�\㊇�#�΁�,��o�q}�3���}x�0M�	�O���n��[���ɺv�yU��>"�B���YhÈ������_	��C�ċ�#sg\�_���Y�L�w��44��%�QV��o�In��j��T�\;6����2�7���ސ��O݂zρE6�wۖU� �������F�=�m�XŐ��Գ^�͸t�$S�VN��o6����D����a�=ϹMJf�|y�0�k�W��;�/�^����T)�����x����#�toESB�.�$���X��A�4��#dɾ��)c���Dcߗ1L7KY#��F�6c��}0��=�=��k���~�����>�s�	�\~�Ϛ!�� �}�O���R��dyQfz���]�'��LW���5�gE}�=����&U$aJK�\��\�K�!�X�&X�����?iI�T.��J��ϒA�űI޹.H����}Vo$���w����o5��,=�W'�+4,�A(�~=ۏ�͢���������߸ʊ���[�^�����]rFs��s��>��t5�2��F�Ks��0>q�,��Q�Eӽ��}]�c��Y{w�"z[8ո�?/�=�����V��piN�# �:x�������b�'�7ƿ}K�G�}^a�2$)��Χv���
���c9��D�jC2�/x��2�Z�ܪ���1��nt�w����OrΧc�9=��oz��E���4$�Z�3$t�w�E\!���M�� ��1uB��ϟ��3zRb=��ʜs��ejR	�3�1ua5s�.�M]:|�|�k"A�+��Y�2*��� �p;ZϚv!��� ��+�q�ݙo���ʯ�ҋ�(���sھ�̴l���<������os�Q�酊/���� Q�UtU�绯�7�Z�+��#[g_��S��ٺ�;�jMr~J����
r�W+�����ޒt�|{��ٖs�أ�:�����1�����k3��eU�d.~�3A�N�ִ���Â̞O�C3�g��q����ГNp�0���'>0��"��ᥒ}4������pâ�!��X3ʱ�2�>1�/�K���4�|b"Z�G��d���7��|Ce��-�U+�N،����{��_�E��~*O�c3���>z6POeM��AU��x��V�OY5Ŵ�z���BH~���2$%����ů8r�ɲG�(*+q�$ܡ��q������E���p�8V:hT��P�~�=,��忦�,��Sy�U�,Ob���aMaP�N~-g���W
���I拷Iʔ��PR�|�cI6kP�nv��;]r�*���z5L�Ny�#2	9+C/j~O���1�4�E�O�֨�v&�*�������潘�x/.f�<=E�N�Ȧƹ����5Z:Q#�턬������/a�'e�i��iOY��Q9�%^�������)��O7�Kxϸ�hqNq^�����n�H�4���5���ϗ)xC@�_�"��R>2z���Z4�A��`SE��Ňg��.khE���͕G^�O|O��60�'^�V���v���$��Ii!� ��v%0�1�W��2��©b1����&�9�<3��S�z�����R*�7�x��ܖn
�bWex��=��U32�\�5�o�W������(2ĕ�}�^��n�։٥�	J��\�
�lno,5��!��z�m�����TA����%Ӗ�
�o�>$퇈d�J�����������9U��cV*�U�������	��WZ1�1�{���C�)�%&��f�n�®g��ӽTPn?�CF'��kEҎ�wFX'�v9n>�i����������MP`-?˅��H�-B>z�.���;C�g��C�~^o����K�7A��|F�%�.͍�>��@���6�9P�D���y��^��(
PW�DM|m8y����-�~�D6���'��@P8E�K��ceޜU��A%���v��/�z���8?������D�N�g�H�����������R��޷�������ߗw��,��p���m���vx�N2�s�M1=Z�j.�J�>z�+>��<�x���:ZQ<|� ��ۄYj���j!�ϙ����u{��`Ǘ�f�b޼�����퍼���;�ʯ�L.Ȭ,Cվ�yժ�ɩ�V�E���c�=�=���;U�-W���K�?�`?��#�P�z�տS�IK-�V����T�c����� �4�"o���!�Rh?oί��tN�٥`YژVf�!e=�N���'�n��KJ��#s<
*>+TÎ�W���e���KS7�~��2�^�\\���Y���U�%���0M0����CdШ/^�����xE��?�������y/r�ŖcrIa��?х���,��
��eX���WϦ���+�<�_��LձX��ޅ����?�Q.��ڿ}�JqԻ��O*�Iȅ9�������`m�M��h0��'b�����G�\ș$��8~�J��*(0vM��y臙��#�K~�0�gKs���m�B�7H�{>�����u?	᭸����f���#��_��\�G�<��˅�s0r�=X:����#3�9T�g0�,e�'�_�H�`(GG �z�f�3b������r#�@yiҥe��]����(�
;r'%W�{�~� %�J��/߹P�R&���^�S{C�V��W���pE�����z�a��m̓��s�f�P`�N�y&���ax�c$6p���ܷ9HCߓ$K��d�K�Z���������Vw�%�>��Y�e� �%��X��ޥ�6���z� ��41߸��݄^����W�,�[~�s��3ٷz�*'��{�8+S�0~�
�Y�FK;ާ)�!��I1{��hM
��q���c��`p3.}�R]4IYf��YK���
��ER.���X�7=�S�J���
m:�~���\�|?H�1  ��%��o-	�DF�Zp�:{�3R\6�L\�f��] =J�=Jrқ7��w�I8��qC�_$�RP@)v��X�������]�^G��$E��<���|��H��b2
��y�}xZ�Ύ0r�nډ��ö��S���r�J��j��: ���\PD��/O�1�F>D��uϒ�������H���]v�
�ݦk�����ң��
����⇡��L%=i�����GA y�t�����n*B����9� ��mc/��6+��f_��������kν�d��' ��b���_��p�^�,zB���\���*�d�c<�D���5�KS�־���4/t�{`�l�8k��ci�(BCv Z�
ɀ_����R��ZL���腀�x��#Z�ׄ[h��h�f����ܿ���rL�:��Rw9���c�[!�lWq2.T�>�j{Rl�ͻ�HP�Z(>�a�i�v�F+���<��r�n��u��5�9v�I,:��1{d��rj��ndj��r�-���o�s�� ��o�v:m���Q�r���nhB��9������5J�{
x�?��E��� �	�:�+W�zד�%��j`��@��YYT��..~�d�qáb���0Q�E�9qԅ}�5��D�y��.Ҹ�#H&�9	%������B4ib�:=Ĝ�ӈ�<����t,�\�Sȵ���xuҼL�۱J�� �R�z���<�3��-	�Eq�������H�ǌ�\SD\��X��7���2X�VQ��x������w-'����R�0�)ڸ$�SkB9��`�A�0�:�����D�]O�.7���S>�X�/P�nC]jn=�����ɵ���ɿ��3X�I�U� 8}�X�v�e7��#@设�+��;19�ۊ��tM꙯�l�i� ��S���,ڀV�*�����jkn>��ي$���xY�2����AE��E\Y���!������f�����j�!��IB��}�u�ލ;�\7����Աw)��rJ�-pf�1C0�1i$��[ik	�������F��	:fS2}e�{��AX,lݙ�����_�]�Ox>���
H��qs����c?�q��x+�9�
)z��ӟ$�?�y���A�F��N��CWɋ�Uy/�է���&��v~�f(
��	g��W���j��3N3X0�G���Dn.�SB�B�?�����M���e���@D	4=���� �({/�x�I4A���~9��>-k~���:�B;���K��5��^�tS�S�`�%*H�;Q���$�<Y��ʙ#?�6��衚�Y��r��^�kE0ךlu�?���ޗ�8�,4�u>͟�������e��@�/��,7���8�2�� ��dLC��V�p}L��X�I u�4�O��ۯ̗��|k�����ЏK���j=�W/�@%��		��<#�&��!�uS�Ŗ���o̊6$���kf�ܐ���|����]�j��$>���!��9n4���b�;�k�+ �s����F�[O,"�eM�@��V���Q�@�R횦�� z�9�'*p��`~��rfL�]ٰ��ռI1����F�+e �
\�w�ڃqN_?���RB��9O&H���ƀ�Ύr�⋔3K�u���Ę�B�&��V���,>Zq���T��駓-�
�C�'*f:�z��x�O}0M��x��U�h� ���D6`ј��O��D$�J�h�9>��aJ���,K��)���x�s��yh�A\s�㉷^E�W���␡6��9�-�^F��2ʋ�<�i)lÈ�����8���!.�f�T�ςe�x��c���F�}[�U�"�Y除�YW�+�t3�G���v��i {9,{ι����o�s�h����!Q1�.KX��1(\�&
?�n���o�<�i����Փ�Jn�ǅ0,7؄�N1W0�u�P
�aP}�����?�KRf��픢���]'rD���j�Z��?֪��k�r���+m&*��Y�� �nf�:L�g����[�}�����h񉷻�#�g�Jd���s����ꇉ�V��[�˪p<A0��o'�����\���g�Y��$�~�*�F&1ut���� o+���jfu;`���ݬQ�������9%{H�<F��6�l�3+wً1_@V�"��r��-0e��{ιx�۔���EJe���cR?S�c�7�]��ʀ#�M���LZH�LE�L���`�A��6&]���ߦ�ʆ�����T��8Yx��xGx�8 ���5����!R�	D�d^� ۞�c���|c����]��K�d\跥���G�]����
�8OX� ��A�k�R�����c��!����U�R�x���h'v��G.��L�C_B��7��0���� ���*����,�P���]�+��w:��s�i��K�S��C�$��rE��^�U*��]�o[��|���Ǵ�*#�����aG�J�'8�岁2�^WӃ�J�����k�eE5zi�U�t�U��*x:	V�#��[���
ڧ�$�0�y
y�ַl]�Xw�V�Q����?�G�:Y<8!��S��m�f�p�� �yDԘAeI���枙�|4�{�P8�x�R���7o�ϳ*zGlF�4��d��虗-:;f[<h���@�|�<~|��Z)��ڤM�Q���"����<�5gU�����\]������ʢ]���Y�g�@k~d��nvveS���]l[���~e@� �4���DVU}a��5��&)�!��`C��	�%�ρ}��g��H{���+���0��+i�B�D�)f��
b���!�!
D���6gw�B�(�R�|���6%.��5����UF���_4X3�&����O������]�Gi����A��d9�vw��r��z_'�g1R����]�1���n���"�:�=F�}���5?i���s��O���l�{���=6.IqV�ٟ@0�:��IT��2�ww/���2=�5J"�c�T�k�Z�����a�A����qZ�Ni����[Y��tI�199��ix�o��7w�U_��\���ѝ7|t4��t:��]�-�}�q�O����3g��봥����/Z=;	q4!I�_�8F1��l�ؘ?���׬��9�l�<������+D��/�+m��ʯč@�>�r�a�^�-����y+<�q�'�'(�cq�:�D�PJa���y�`�r�����s�i���,�S-k��X����{*\�.?�}G@�RAOe��g���d���A��)�BZ�*};��V&���R��؈l>���x����˞D Z�m�C�Wy��\�Z�\�Z�^}6U�N5�����wp�uPa{�:<���g{��;q��	0��?��Z�AlO��=D��)?MS���LR{�~mB�����@���L�����d�v� ��A����S����I�Ei:��W2�β��姰7y�/�� f�ݡ�i*Y|h�"��]�� ���۪w������5<�^��|�]��sύI��,S"�y�HZ��,z��D�պk��y�]���!��L�jZ5���J*�&/� #0:�g6w'�wy&�ѓb��5�7sy��8�u5!�v���K�����u�'��J�2�������҂��7>.8f|�Ͽ�s;��m����W��@+:`��k�~�lX�L�і��჈U��ҥb��2�M/��i�㓕��͸��%����T)�fmUsCy��jmk�TA�4+x~���e--U��<�l�4�O�u�����b�廔�A:��rd�[$ة�ؕ[�2�r���hta�g<7i9q��T��Z���h[�]���=M�Uv6���2fha�HE�M��y�M9ޔ��_.D���8Uj�w����O�&A�� j���9��ު���n-Ҷ"Ezk���N|�p)��$�rnW�E�|3���~�w��U��MY	C�9�_n�9�[�X�J���|>g�.V�Z%��6"�6�s�EׅU�w��$jq�,�t:� ��8��1q<.�jд�jh�n6���&��l���(��8�9����8���u����̬�L���L?������U^��ټ���DD�����K�5�*>Z�vuf՜��W��E��4Ld������|��M?�f|^�AB�_6���9F=,$�=h��m�H��RVMt��54�\��_���.���'L-2/���͙bUf!�/���ȅ*��#_~�& �0t�(�����7@Q�wK�#IW�a���׿�n�v�ru�}LD�o���)Skw0����!:���I�Pm�Y�x�̹�v.H@����[X����+�vi�;��E��v��=���Ɏ�u��ۉ�u���&qrɊ�@�v�=�a��jhͅ�RmZ�e���}οó��Y=h?ߜ� ��"hU��3E�*2��"��|ҰC'����YR�d8��ޟ8��C�U�u,��?��M���k��^����P,i���Yu����S���Nf��4.�zS�,���N��m�Y D�,̇���s��� �E��A�P'ZlZ��I0�������\Ȅ(��d�X�z#�Ͱ���ĿŽ`4Y����#E���{55�R��zY���[�J➿@�Nv;�Ԑ�y[���~��.>�,`��D�UUԸ�ǬէO�1ԇ�<�d�ݕ��\�q�����T�XEO ������DW�.co�wֱ�yJ?�;s���*ѯ/r��T���Ͼ�����X��<D�@�J�T	5�M��H=��i�Ȋ�_]F�'+9M�$�x��UUk�Մ�\���ߥ���/�	 i�����p�]i�S��z�n��+�0/c�W{��e��n�	Q�ꋔ�낥W�����nM����g����BO�,��ή���iM���&�z���:VcS�+߆7�N��}�
�Mg70]�-�ﷺ{�X��2b�̢��I:�Ĝ�}��Fi���¸��װN8u�oT�W���_8��lH�׵9!�?������DGZ��o��g��7��i! �@o�Z��%�\�ʻG:�EhH�Hl&�6!����=P�0$�˷O�\�+�q򈦘<�uSLC%�E�����F9U�@'�1w�q)~z+���7x̥���k��vאU#&���${����ⓛ�|�i$���SG��7�v.�p����q��Xk*��c�$�O̝�ٲ����Q��-�By{���_t2}]^�7��	ߚz��_\j��=j݈�#�������Niq��V�������ס ���]$���B�k��P�(���6<��p�����>	[p�-u��d��nn���݋������W��R��#=ཌ��S4K��"�v��E�^A��f�
��m�X�4�W/ h������;����� ܤ�t����6��/�	&����/J�R��wi�j�����9��!�ꘈ�'E�)��"_�?�����!$*x���bN{2���V�ur�&�C#>y�r����,+�0���E���;��~��]����ϔZ�.� r���|���"��L�5��WL���5>��,|���4=�tY�~����Ö���Y���7�W�ߖ�V�����]�F::�bL����nށƥ���v���n7�'d�1�F��"Q�$X���,rp��}a�$B��e�����
��+�T{�X�q`!Q] 斦���]�����,c*O�N�сϚd��g���H��҉}�*Y����̌�ѣӮB�xC��MV��&
�l�
����K�I�U�?t�]nP���J��AR\Do�qf�xp�q5x�d�k^� m"��q���zZ'�w��[o�m�*���o�Q�q~���2����y ���@������	d��m���.z�G'Rp��O�-������	h���&�}�� 0��%I�	�j�&#���sN�=�X,s��i .�)"㗇�7����%�(��i�e�Eg"9TFA��E����=��l��U��6��Q���5R���K���N��>��a��d��6����|g�i���v苧�i���*�g�L	�g'��`�~l�)s�|<|�o�۫��,���8/�v�@9����#�ΈЏ�@�~�q�ǰY�i��̉ZN_��Kc{�	���˼�S��B�؁��:[�?R@��Iyr66<�΀���H4��P#^8@��x��|}�̌g�����T~)�:���s����;�D�b�O�m-$�=�>,��r��Z�玪�a+Z�瘠'7*�S�[�H~%j�o��}r�+�°)��:�r���hx�)_�2������U��l�a����y�%��aO�b��Y3��
����x��y�� �4V��2�cj������(Dˋ�?�f����g��Y$�:��eWߑ�~���i��_��W5ե]�*IX~�9���-ڤ��0�^�[�`P���L�l��G�]����L֧)�Iqr����L ��)2}��c��!�&ʵ�]�����-Z�z뺻���ؒ��U�eT��-��pݱhpC�B�o)�+�W��[��-��3�?*i_X��\>VnTs��_  ���+) ����t��°<��k����p��l|�~�D��C͖[�  vz#��ed�]M�a`e�jD�p��뇩j��2�a�Vq���6b�PL�s4���7o�@wh�ȷ*[��G%�u�#����.	=�}J�XU"�ov��ā$��[)g��TQ�X܊��:d���ѠV��X�Msar䃽'C'Ƭꦺ6<��A%���-s��	�Y��a����ؙN{��E���O�4�ܧ1Y�p9�c�u�%�R�|��&�զ���W��׽�E﮼��(���	�2�������yft�!��3�G�mW*����ߔ�TU������~���c��|`��N�����5Sl�_JL�wm�Xf����lkk3-q�[a������8���I�� �#�G��)����h��C�DY<�?I�V]��ٻ{6���9V7����$����{�]L�&]fJ�hψj��Je=�V��A��v�4W#*����uP!����V(V�zm>���G�ؽQ(Tm�enS�5�,���hyg��zd!A˟���շ����$1I��@��ė�Y�����Fh*��$=D�bg����̞�4b*�#�J�Q_pK@�5�[K�vhf��O���'R�F���@����|b��X.���6��L�y���a�^^�/^���0�J��ʛ�"��itO��$�o6��% ��gv�x�-�Q��&ʔ�(����b#�/'��CTҝ�֎�+����u�߇��3��w��O��>�B�D	�����wB��=v�萾�3�Σfs��Kl�V(,� ����门�qu��1t�1�ux�*{��5��X�B�p�h����5�����0#���/���ԫD��?{;���\�R���W	��;�m�/�
��[-'+K��=)(�C�G�r~��]���_3v�U�1YQ��*���:ni\֟U��מv��j��]	C�j���.���~��j�K)����/�P���'��C��{f���wYШ� �=���]����UV�F�����!������eO��4n�.�<�{�O�[���D+��j�iO{I����0��p��U��_I[}=��4��dWu�8�V����t�O�+��%���KU��<0}P	��X���Bf�Z�n����L��)4�K[�`��3m��
�eȂ�e�
sH� V�}�B�/�M���{��!�*ꆬa��zb�"7�q��'�n,%�ڬՠ|%x��SJ~wu��mvA�8��)�N�@����:JJL�\�O����T�E@���2q���O!���&9`�6-.E�6s���}��3�6�1�8��d`[� 7[�s�n��	{N�'aT�;:.���:�+�*��yF �h/ԓ"�;S�}�?�2Y������L�o��bC�3b�˴�sV���=&YU��=��8�_��q�)b�z����z\(a�'M��D�.�"}ݫ�w�����`|E��P�\f�6 �&�%�o����?_�~��,tI��W��jm�8~�픍��ջ��@��OV4/D���\ ��Ehv�]��*H��P�!�^�¸��Eoa��&��?�xC$��WV�͹�r� �),�?WsY��#��]�v�&��ļG�F�X�\!�Nl�R�w0r���Uh}�����O��tzz�,�!��c�/�լ�8�%�ކ$�L�G�)���}A-w@&���7�Ȧ�l����٫Հ��?��������h�Gӆ\����?b���+_Mj��@6fǬ�a�$�Po�#���d�ݲ)��/��l�ɝ�O1]}ZN�ZV�1{}�`w_;�ߦ-�,�̨��iw�NF�o�~�l��R{��D���H��̭"��uX�ҫ�ЛFװ0<H��ȶ�]>z�
���j��2�ۨ�y%�u��R��¤�<��R><�A?z� ��ߢ��r�u�b`�;��B04�I�A�+��a��'���3��y �ֵ�-��Ū��Q��(6�qz�][�*�����\����{�k����>!������]\I���r��MJ������tN�h��x���b�4�+�FKx�S��,%�M�_�1vm�]
++��]޻���"�#�O�sC���U�U���b��i��<�v���b�+�N�>��a�K��ij��N��z�dg��f*������?BFy<� ���m�I��@k#1����P{*���R�����e
z�˾,W�Z�G���>��9��򾠏�b�5�a��o���G���Q�);�f�\�"eu)Ucˣ����ن}%�|�6��}�L�)|23]Up���i�2_�uU��k�&G�) �D���F��=�|�>M�k&�P}�YXE������.�CӯsoO!}�u�-�c�����1c�����5�"��*���@��޹����A�}���]������\v�����9��N�i�֩*L��p� RH@`i���!).bn5y��w샹W3��7�9c$XPw�o2C\�MI�]g��PX��0e�:J7[�x�,��,C.��6�\ґe����مAʄ`��^I�6�{��l� ����	��ȝ��߫n��ڍy6��D ��+6GC�S-�'����^��G� �p)��M�[���)�BJ���n	|�~�.��t՗�j�qm��)�>hSd�� �4��رQ���i�8��ɉ0�+_/%��22��O�b:���I��7���Q%�/h^��u�(Eζm��٥���O�˶x(=~��x�tY���.������������'~}׋ ;�U�g7�K����P0��3�Xߛ|w���gh�L����ď�#!�t����Qt�O��������1��Ha%^�o��f��g�l�y���(Q�b��/����������\��x�A��;`����>1ː���>�,}�1�t���Z{��뗕��yj4��&����TJ�1N�^�-�I� �ׁ��)��#
�����r���� �Q���ӂK���eb�� ��  0����x���̞��?����=i�t�mڠ{�֦�E���TC?(Z���j�S���P-�7vC~Q}��6���-T��N,�O�_R���.�8���xO��Y� �W�W���L�@��A��j<�ā�V�P���F�1P����P9�s�z�j��n�vé���g}�F�;_У�QD�^~��S��څ2���o�O���1G)ڛ>����ȭxO�X�<:�hz2:���]K<6?���A5���������D��D� � t�!l�{"wk]3������f��w�#�sr��̾��m���M�H��%�cZ1+�7�X����g��D�����h�L��1���!X���t������ ɯHEa)���-����B{�E��m��F�����o �SB�5e���o��[��o|Ȭ�I	vf˃���cc��A!U(�p�^��@�Ö��C�t'5����Q3�U�۽c���G��e~�&ml�Qpsb����J�hf$n��Z�L͵�f������Owa�?������0l;�}��L��b�O�����%�{�
TN˙#����(�<�?r�]�LU]m��40�k�1NY�/?n��j1<H���jQ�s=�u{!�>D;e9/az��L�,Hn��މ	�,�ns�^�޲��mÕ��yEhD/��H��@i@`�G�$n"���ښj�ѹ�@�<dzI'�0��"0�i�/A�0��|a�7��#<�6A#���>
�K��a�p���S,�H��m��,��bA��� e�y5ڪa)�\?`�ڤV{zx,a���[{�ɤ�������bv���Gg�MĘ�̋�����ۄȑ���ꎼݪ�l��Z��c$��ݱ�֧m���Z,b�����sx�[��̯V� �;�5װA�M�Û%�Fd�A�����NA�H���8�g
����bqnN�� ؂��rT�B�O�(�z1*=�y6�80��}p;S#�=���B/�@1�+���d���"K�f���Sҿo\~8�HK��g�sv��d-}2����@�|y�N��'��E44�l���?c�����K $2^ nwj�����/��x��r�~6�!�`y=�̀�?l *_�_3΃�__����(>�6gVU\�K��2a �3�j�e?�i�����`6��'�x�6�r6+���EW�o�d����j�$�4D�2S�[����|f� .���7�2*�Vt�쟽%�e��@���6 
g]�9
]J��������q�a��NM�����Ksﬔxj�c�Ŀ�+Z��ڀ�W���;e1�4�S�K�K�-��9y��w8l�s�4m�YnP��}	��^l�j���fS����Z�Mj6�3�0�j;��bY��wL� ����NB������\��:�:��#]�m����@�l�9*ө�\s՟W��Q�#�S7�G�n�s4�� 4|:�����hmd���")�fo�D��?goO��p"6�V#���}��Х0@z�Ϥ�{'�������U�.�S�vw���[)�7ܟ���������5_�NNjGW�:�����S�Z�0�m�odE���˹�t�G�����kx롲�i�d��V**/S}��p���Ҋ�Mz/��N�f��a�T�tb�M�}�0?bfBy���!\֞҃�r�~DA�N|Ed�vE��~��PY�i��_����;�f�U�k��,^D`(i�[i�O��G2%�Wy��y�P���Q���{��	2;�!z�����7:�/.Ø3�8��_��)��EZ�S3���hVt&���}z��O^���E.L������:�Q{��ѵ(��yD:ʓAtf��g���DZY�%#.Q��;�#��ZnnzC:�����&E��,@� "�O�~[�Y�d��\or=q�:~�S�#�U����5�4/2'T�_�33��5�$L�m�\��.y�z�=sx��No�D6� F��%aX4����}ޡ���P<]Iz?]��`�s�;n���H@�v����omC�	��ɘ�q�R'�d��Y�O7�����"0ŹC܂&%C��l�@��]���	^�$�S�q�[���p^M�`�}��K���B���^�� ,��SE���}��VP�*�Z�R�LKC��;/�'�}��ku����__k��n��12�����%;�N�����w�`�P\��gKǮ����'S�`F��$��;��P�\�=
�F�F+�z,������@Q���{�`T�L���?XĻ=��p$�Kٕ�}p���6�=˯�������4�h��Jx�'?H�=�q�5�%ΐ�)5�HF�з��|�@���L������"��p��^+��U��@[]ƙ%�Ot(1��Hz;�x_l�#R�m5x\"���(���X��Y��y"�3ۀ���/6.�����5�I�u�h��!�)^��ڙ��!R���ys� Z���]�xң1�:�,�CH� נ"��q�K��T��
��!{�L6C�����69�~���^����+��.��?�e����tTϐq[C�m�3}��vβzʐߏ}z� g�^=��r���I)S��鬮,D)��Y�)-{ʌ�~��1B��:��t��Zޖ���{.��ݱ�11|�X�6
tO��@�_��ۯ@�r�kИ�s��/���!:� T+b'����_�whs�}�!h��R����$?h�{eR�b4�Fd'�����r�C`/hМ"�v�%ғ�
�:���m?��d��&�`���%a?�}�Un�9�o����߉?r9i.����m�\qρx�:�VM߾I� :}]x,�ZV�H;�e��,����X n�
.��ͼGH~�-�k��y��*}��k{�i��ˮ�AJ)p\��7��[����Ҥ��� ��N���Ӆ��y:���[�m�wCX]���B��.�=#��͢��J|��Қ!Y�^���&\�k
��-��X^BZ��+(�`�m�E;��G�
��c��S����I��FDۓ���z��;�0��_���.O�Z;#���9�5�0I"|��|�b������8�lޢE)��r/�7�|b�o����,y����3�b�f��q�' 9���i���y	��XKc����(^�#���y���&��|h�X(��q���	�/X��(:S� �<+m*<h�?n�Z�����r�7�a�]XN��t�EC�2�@O�����֤�?����<l`�t�=v�}�����e��)��F������p#\����ܮYQt��Z`�`�m~��ψy��Rz����S�к����.f�7
�Q+� �
�Ƨ*��ð���^0n�pJw0��e+���	�M�&�;�\�Ε�ܒ�y;���^�_��:=�K�#@��<����)h���i�r
o�~�C�6ϩ��`x��(}F���@l�e�eq*j)����h�yk��)%l�͓�}��t6�<�Y]
�nZ-��}�Y-�i�6FQy�X�����8vmq�&��v��8e����`��.$�����.&��ZM3(��a�C�>9Ȑ��E2H.7����L��#������`�_�)���m{��pw����p��;����V
��T�5���}�C~B�,��&`)������S���v���T(���sN\Q}k�@e����Ǐ��̑g�vԱ8��QtF�#�H�`��n&�g�:���pG�ԑk��͋��zR͝�T��7�N���W�vAB�?��-��H�Tjq.�Lϼ��_߹��6�"����oA�lx�]4�H"9Y[c�}�c��ボ�P�h���2r�h�����M�׽ǅC�����q��/�fzV���GS��Hۈ?���9>c�u�*�y�@4`��~X-5���f���8�w���Ķ�vL�k�OA�w�f9<;��+{�m,�� q9���'-\�۴�1w�T�NtGߜ�@���=�;��ifpϿ=��s�����^	D�S�a'33C/3���F��,%*��^ƚ�%�Q���[��K{�fI�'�ؙ�^!�[3�T]O�@%�F��%;ٝ���)���"���냞��]A��w>jU��N���v��~vI���L�،������Tg�7�����#+SP�Vd�:�=0wL,�̬Q]��;�50���d�p��H#-�������R�ک]�RZ�.jf.�H$鱱>��-A��G|m���Z�;�-:Cf���%�np5�3@��jA;����oO�m�*NgY�(�F�^
�9�����s�$�
�#e[�?��Ra���Y<vsB�L�}��W^F(I����?�%E���D4��,y����SV��?���\q���'�� ���e��v��@2|d"�p�ccS������zjjj�,��K%W��k7�Ϗ��ֳ����2۞��u�D0*Jl]x߂��ơt1� ��ڟVې�-��7�������?��ܨ2�4�ɋ��hd�̋N9.S-�nr!�ӹ-i����i:)%�	ʰ���M�
y�lݼ<:�<P!���ڗE�~g�O�k]FM��dۨrq;��gZ�F)��
���ڲ#��}cv�s�N�XǤ^��ɥ0�'(��(�����JY*ju-r?�U������I|�]��"9Sxc̐%Y�����
�rI���'Jto#�n<o.��y8O���b��}%�X�����$0��߫,Gb����
q��c�I=���`*tO��&�	�X��K�ֻ�a�{�u��Tc[X� ��m�G�S��n_l��_a�$�V>�.se)ӊ,�6/��ՉX#�u_�_W�q{��pf�zƚ̊r�ԟ�=��>�9��y�3=}��t7ͣS
�'����"�L���w�pb���UɅ\��Dכ��(ăD��k
�k��-D �_�YG�:��4L�����l�ۯ���]�e�;��Uz�S����'+�!b_�ԭ+P�{pY=W�j�ꖮ�������R[��tO��7vJ�ͭO�$����^�u.�3?^:�mě)[?�>������$�o|g˽ݒ=���j0P���q��
��4;n#~�h%���2([�Zw�w�G�����^�K�R�%:t��gW�4���O��O}MMf���-X���YE����%ڬ�J��;�=\[n<Y�
�1���<���-wp7ï����K�=xw�s0E���G��[�_�ty@�5�{[2��M륀�}Ѷp����K�@�����fU�].���]/%��RK%��N44�ͅw�sv6��[��C�>��BݼׅL����������;)Pi55�$k#���I.�&�wY.�=�� ^Y\�K: �\�u�
O�lƾ��ܝ�|�C>��4���j����Xo�	t�<f`wC�m*�� z�7;ڻ��2�D���)��`6O�R�L�*j������8M�����u���ڲ_}�V�\�?q�{ӗ�M�V��J�J�t�5�4/��E-�mEJ�X�<��|�ŭ�j�"L� w?�rH+��s��[W�=��38._?#9oI���a
9�s�j�k�Η�!�g�{F�f?�O�����>�́��
�ܷ�|*&C�� <0�Y�˹ŗ�~��\�{����*�/�ᶃ��?�l�;Ky�8B�i6��i'�~<'����_�{P�'���t��%������S<��'~��ƨ���w�+�S�mCI�M�o� �����R���m*Sp����@Mf�h��kAE�.��� ҄`�AAP��K﨔 !eW#iJD�F��"UzU�5���~_��yo޼;���3��9�w~����c�uxߡ����ޡ����{�@���j�,G6_A�}H��\�8x�T�ǰ�G�umn?�8�ʽ�Xy<�5�߶RZ��Ri|k�����BV�]\�0&
�#pi�/���|?Dq�b�/��H`J���j3*� G�]�q��0��Y�
��5F�ֆ��:��W@�Z����[����""���H\�Y�T��H�`������t�6&4\�u�3�3b ��z奋�l�g8t�~�{C�V'
 ��m�O'C����t��J�nYS����] ^"�q)�4�H~ e�@ޡI�+�� E*BY��,�D��	W�;����1���]Ǭ�w���F����ڿ�?���m0(�-�C!�bh�X�t�2� r�5EYa ��ß�,K�����`�+����� �"�ҨT�Y�X��c�Ӷ�;�����,t��i��C����޳`��!��w��iJ�H�n���yx�[����C�@�n�>����g�|t�b��D\�^�I=�d
�Ko �PT\�
(0+NQ�1f7L�QF`��D�R���޷A�ؾ���a���?��!�8�u[2MX�T2s���d���`����D��%%��5k!�M�Ï sM�z}FR��̕��eǵ|��C��i��ل��(�W=f9�:�U�) ��V��^>^Ul�V�8_�[>b�hY)���C$�2o|���|t;\�W��t�\'�qb�Z
��w���P�� ��-�h���Z��R���t��Y	Oˌ��9���d>=�˹�"G0�����7�c�\}K,M������*̽Q�R8��v�EE{�Z�Fnk�)���ݼ�S�gH�S���&ӝŚ�^�n�v�����CX�|�N��A���*q�����*�Jj��^R{�čY��㍟�f�m���n\�?��y�(�d��Q�i�g��i�9��;��=ʍ�j���Ȟ Y�y	���qz�,$sH"�x�)��ܷǩF2�A؊�j�v�E���e�CD;���某�h%�vr��F7�ފ=G���&zO�����|�V�(E��1��*�`�[6��>��a���^a)�E�y�g��K��)������.�^�l�*���Z���䌛���������ʒ��3|�+�>oo������w������%�N$5�$��]�L ��E���-
%�*�S��� ׉6�OÇs��YB���Uѳ�-��'��A9|��KZ�Z�׿u��]�
%�7�������9J���[�zv<��	S�Ǆ�ߣ��ĘAN1�[��̨��A��\ۙ�������*�w7I��~wj鶙�E�fnoظ�X������XǯVә��u�U������f�����^�S~�4��O@�H��7W�#PM6�J��^@�k�N�Ǝ���,G�Z<�?��=v�~F�{����Qk�n�{lw�mxU�g�\?ˏ���۝�NZOK���S�;�`�b,܂/�q!d���Y�4-���$�ob����b�63V��K��{�փ&C	$ww�������s2�Z� �}l?B��?�n�=lZ��F��r%;?@o����[̰q3k����@���V�|Sr� :��5Q��@�#P���D*'���m�ƾ�)e�b^�wj	ZE���B�6�8���פK�9���R#v� �����cK���[�f/��>"���L����z-��#gn�6)8B�8��2D<����X�����~9h��;�d9�Ŷ��<�x`sʵ]n��f`1ҪL����\.V�YI0�w�]h�k9���i�A��3�ٽ8@�c7>��oח+���H Ԑ�aO���Kf��)�k5�$û���V�egb���y(DX32pTw�a�܅-N���o�J�<��ݐ06y��
��}1�v$�o�&Y��+�;�Ln��p��Ţ!3	Q���3M8֡1��b�Ӑ�J�i�B��g��ѻ_������{����m�t��XG���]��th�Y���&��k� ��҇�O�K����{<a�L��۟'�¼�S�ma��e�5D���]\�?}��z�`d�֭!r�q{�/�+A� 	@ (b������SD��cT�+A5R�w$��ڼ-���"7��ɱ��<��(&�>�?O����T5B�膎P�;� 1����#@��[Q�4{��Zh����C�mf�_��_�=.���2�(Y������~���/M����q���C�6o���ţ
I� �]�=�	zy�Rѩ((;Ϧ���w�o���p�{���u�\�\\���M�0�j����#3Y����.���[Y��u�u@�ƕ^��A���I�#�S���D�l��ǧ�PG?u1Ì���c�[Ua�2�����������Zr9��!��Q�u:\o@�,�s�>�ƴ@�_�0<R�v>��Ḷ�)���ńK�:�y�xs�H���v׀�W� �C]�K�%�dm3cg�ou�(<�_���,���PBaᅭ�H">�X�#ʧ�lQ��j@$��hc�rv�=-"���g��t��IDy��s\n���` �M=f?���F9gsDMa��ݵ�9�8_C|����l��'�9�pn���+���+��)J�:��ryO�1GIXUл`�QH�5F�&P�T��>`"
d(�u��A��#�,Z�}��m�:���i~U)���?<$x+6���~��ԘG�q��b(��*��KhmzX�<Uz?�S%�(���r<�v�k�=?�i��=�T�����V�����O�d%��HL8*=���� 9hy��+�0^�X��M%_~�G;��.^Ґ���?y�VKy��@zL�xL_^�cw!k�A��Ϙ]z����&���]�K�[5W�uc�ki���C�<����y�����X�NEi�#�.j��|���v���V���Mʏ*��f������wt��`���Z��^cT���Q�����S�Ǽ$vl9���E�g��#Ϩm˶�\86�z�=�D��X0OM�̀R{���{%��U���-c�8i����L΃��JSӂq-���h)pM֦�ƿ���M�oms�;+|��X�a����'��hxgQ�\9�]�� 'TʼS�d`�����7�;��*�3g�.4KN�<��p�Ja�RHF�?�6�7U7vV�������mSbV�V*�㇃��OOM�h�� ��"/�Cg[*�}���=w�\;���B�uJGuYC�	��Zh�Q-_��q�������"m?j�o�Ցjm��ӝ?��㾋V� ] l;�1��
7[3�I
TKk%N��Fn�X����G��脝{0�U �R@�矸~�.7���lՓS���K�ns������*lpoO͑�Z����G���Tk�AM�&{��v���M3p��Å�ǂZ���v��+��WF��震4�	z�� �A���
��ng܃��P��ҍ�٥q��<_R��>%�ր��$�(�$��p9?ɯ�����-r��3�`�JQ5R<듩���	0����A��Q��^��r����&��U0���!Ӑ<��������|�Q�������旹�>�j(1��+K�~���<��K~��SO���p���/f�����I8�����͡�"����; �:[�]yX�������9K�q
x��u뎨�9�P ����[@��n�Y�@�P��q�KRpQ����%����z_' �#�~�Ti& �����M���Zz��L6��?O+C��mG�g��TB	��8��}Ѭ�.��ƾ5�յ�$�/���)���������ު���dzoΡٲ�i����Z�Rv_�����эDT�}	�%#tyVcA�,x���ٍ	��<��0��(�pz��L����d�b�B��'?��F��Ò��ҭ��׍���s�7&S�C�ƀ�0��z&�4��cGδ �������ߒ>���Һ)�<���������q����U��$�����圷>ǩ+qK���um�;#��K	���?�zN�b�|�Xn���QrW��ax*�ކ`�p��.��Yn_���%�|UeU�ij̵E�(8=N���q�Co��u����J|S�I���L�����7b�B�4��v���D:)gy%�js�m���29]�@��U�x�鯅�����k�LzƷ��{*�9C�s�k�[ ����Ť��n�s�վ��<�{��*��򍛤���uu����9��& �nuЬ��|$�_ l5��c"]���ZT����:6��4e��M�+u�!p!y兖�ܦ#��O�{��Amt��*�yQ{In����@�^�4JN��,�T����ު�j���Z�� џ��q�DZ���+�)��"�v}XyD[g���]!�v���7r0����Cܭ�"��;�ծf>��P5 �O9��R��M��G�s��pY�>My�gL0���ƷS[�q�H�Є�,P�\mT�7w�C�E��:�`EBr;��a��N_�|��,�9ReI�Z���I�Ifn<F���.7�I�ۧcꮛ�3۬�̫�T3�C��P,���ؕYt��᚛x�T�J'�lW���tv����ZE3{˽��Ty�	���,��M�n�k���l9\'g#�gJ�.ׅim�`�+�A�z߱�^Nu�Yz9$��Pw�M�b�w�d�ne�T#�m,���:��-�	(�ʚЎF��]��H/�i����@>c׆�ޟK�Zz\vm���3t�o�E��Ƌ�z]��C)�F�,:�Ұ���~���q��	��T�ۆ�j�ə�E�ȝU���)Xh��v#W��!m�wb��E�<'�DQi�o���+CCI�=�B�Л�&U�i:�2x�\Y"DA(z�Nf�$u�	ښ	��������: �l�Q�<ڞ�\3��0�|~����ZռY����ɍ���VT�ϵ�~~�Ck���K������=�7��&�`�E�3C(k;
 ���=����3���+r�m�T��]�3`�tj�������~^��̷���y7xMZi;�+�C�eA�W��i����r{�#I\}X��{ɜԇ�X� �G���c��}DV����Da����6�^�a溺*��o���Ǥ*�tv��9J�͗�f���e���«�	lM�.���u�آ6�[6jༀW���RSX���[&ݚU�dA�uBɥ$<�
��2���V�����$��|0y��j��
���.lZ&�I��[z��<�fO˙z�[}�I9�ܳo���'�w�'��Öc�����m�t;ס3C����i͖r��΢2]D���!P�	�����o�Ik���B�ˊ#��߲
g�7�r��Q"�՜'����4/rڋ�����4�
xx�RZm7�6���]�p��I�7w�6�rO�#��[�ZC\<�[��bs�@��,o�`=|��B�~�
Ji�Ra�@�܄�w�zf�,x��k�ly\+���o�ʨ��>W�^D���������7ŵ۫8ԅ�r-�bl����b��uE�z�9�F3��c�[���p�t{|e�}/��E�HIϳ�)I��ߞ+{��۝�IY8z��w�`���7Pi#���ћ�]q����fX���'�~��eRnW��b��2��@�U�{{�#ZBT��ـ�􄀨{~2:��uq{!$��h:���D5��6"�,�T��T�]�OO��X�F5&����yc$�����}�[W&f<~��+?W�?��K¸�n�����B�}��O��k�.כu�%��ĸ�?_E:�;�(�� �/����2����N�J�)^�6�/����F�Kwr���Q���*G6�����Q��g�dE gf��l�X�j������sm��)����n��_Vؽ��^e��p���>9�J���s�����gs��`���&�`lS����/�8�mV�b��_c�E�xd��Mgg@�@**�����;	��_����"z�V�h	�
��9�ă��;�T"0[xי	�����Aw?�g>bT���~��/�}~����;߱wˁf�\oSS��_�zU��� /�@>��יc�C���H�U�kB�^co�<�AE�Y��'�Λ��,�z�ri�H������C�6/���D�̻?��_1�F�dz�-,� ��P��*��������M���c�^K���L���^6 T-um�JF�F�w�}�4oI�����u��b�����h��ӡ��]vlMU�vou'����2����rY =uLa�戄q���W��������!�(H(�<���A�GB;b�� ����	�)�'�c�7�����)�����&����6�6�	�x>���^�؟ն��sH������E��]&� �����y��=��;�5��_��d^�N�ߎ�_�8Y�1���#�j�i��/S ?+Ӿ���&�⮖JΒH�,��T
�����?�C;_�(��,��B51�����h񸊘�c�nr��<�O&ƭ	��3�J*�� �E����-���zYP�ԋv�m�N'�tr�L�-��<j��n��v���$�mz���0V{f��k	D�-�m��c����E�B �:Ɍ�7��K'���KC!&#������?�d����AЇ�3`�~"��h/���*r����z1�1�TWo�hj��g�t���(pg5�p�bY�7��խ|<!�E����jb��j1��;zbt�&��"r�3|�33EBoݺLZ6*���gl@�&�g�i�{�V�#�s���`��N�u.q�Y��2C��S� �*�g�s{^02:;�h&�`k�/�r��'���#�>�2�#e�;��w"�s�Y�� d�2�`3�q8c�@U7�y@3py��8�$˭��h�!�A�Q�S�-7~�I�}�����B�B�}�����\J�����%ʻ�)�y����E9�&�{���p���ĵ�c��� s3�c�p�Á��q���R�R9c�Z�����+�
�vQt@�'u��$�B_Q��2O�h��ԟf�ɞ���z��W7�h��~�����j?��H�d���m����!�J="��Z�� :)0���7�l;�0��@�
�p�e�_ ȟ(I$�{]jmrI�M��L"\�Ǉ\��3v* ?vy"9�=Ma�y�������c�e�D~KcG��#f/P+�^H�h� �_ڼ�O����p��b��!�m�<x�+���un��fG��ˋ�7�-��X~�hc1هB���~���.���E��c�p��f��9��^���Xu�:3�E
pF�{��p�ߥ�YA"�����.��uk���-[SGZ�6��3�h�*��������6�WbX %� ���[l��-�&Z���QZ.3�`�iUN���w�I�^��X�X���|w���AE�s�K���i�3�K��k��d��K�J���bKH���c/���W�
'߇������쟇BM���y�πެ�r�5�X���	�:��2������?D��ʕ�*��5R݉��Y �F�}��7gLj?�$�\^��4�)��9d�w[_b`s ��~aRk��(�|��S�%�0s6������C�;�t��������|Mh��B�-7Px��C�vY�@\ה($��J�e[��S)����~R廨ʧ�"���]�c	������'S�F��H���7N���G�x��Esk-��![�|�Y�8�n)hTY���{>�ak4��G�`�)���F&�l^NW|�S�J��> �%1$l=I�M�h\��ˈM�a���
��S�B@�PgC)��Nd����-I8㼔��D�:�v��Er��V��-_�h�V ����﬘�%��@��ڨ([r�p6�5�mr���MR�����R������sz^!#U�������`��a�~�XV��T'�`yz��G���^�
�j';:��8�=S�o,E�r��-̔:�������<��'�]���&���b�,Ԃ%W�+h�U#)��cf��V#Z|<�t�Ư������Ϭ'���+)p�4/l롻��j������c��W7V��Qo��ۢF�c�2r�`Q�/�f���L�s��r�q����~�h2LVUY	K�j�f�Ne�ƚ ���zFi�o�zV�N^?�+�$���J䴾B�^G;�0��t��T@A?{�9�� 쿸X��>�Rl��Z��4+ǿ6{]��pD����'d�.�5���3ڱ�j}|�\��n�ys�8v��V�� Z��8���e&���pp�Em���'��_�A�+�c�NO�F�Tȍ����*&G�����C�頾QN�	+z��--��F'���D��7M�v��6^Cz�Wl<��Z*���8m�O��y�K�g/���
�?�S7{� y�;#�Ժ׸�p⁨��_����O��{�,�S/�5{��8j-O��5��ӡ1�^��P��;ݍ��g��>�1}��1��J�Xt�7`?�x�o����4FD�qg�	�O=��i���`?a�QV�y_|QC�Eջ�Vv�u�^P�鹲z7Crd�2���񈪛�}���w�y���� (��60��[`m�yW�������ms�ػ��4�~I-��=���3x��*<1�٬P�n"Ǡ�ݳ��%[nW7	-����l(�a�t��,�H��V��35%�EàFa����..�vD��Q�I�LKn����"�}'����T����f ��0��%�>�oz[Ɨ���\����j������g4m�Q#�&g��f�L��)-[��d@$,_��z{D�J��v	`����{�����Ȗ��� xY��f"͝�6K$�\D���u5c�f}	�P:�mQ��Z�j6�_30�ӡ∕�u��TZ�ַT����
P��ע��%Vq�����߱������[��
*�����=�3�R��NK�}�^�h��W� �]��m^ќ?���Z����\�V�R�Z�s�-��!��l�X>(Lֱ8�DLDc�T�P�.�a�<�f��INn�!�D_�l�[��[ AU��|����Pn/�:���H�����/�N�#;�E��F�d��|	�@�����h��Z2K�^��T���R4�Y	n���]/�?���r`��[��<��Ht�q6��o���%	�^�2cj��捈�+y ��*1�,��Ъe�V(�K��j����&Y�T��B�8ȧ0ק&�[�Z\p^PQD�9��Ŗ�M���/�lz9�v ���L�<�t��#�LI�B��5���!T��t*�BڹR�R���#�h��kZ��k��#OK�yN��Y A��/{��� �S�X���)�ﹷ��ܬ�o*���"Of ��k���
�6�n��8}Iy�(�^����C��D�;<�>��I^@��i`���$�5���OxnL�z
H��o12��� �&B��c��Vf�9��{V�T�w�^-A8y���^���8�բ��ia�
��������Xօnw�]L�t��Mj�U����8�G��r�bX'>�������7�q ������I3gE*4�M�2;w�U�uC�y���}���3��qy�Z����&�Iݮ8��]4Xx$J�l���S�Z^�q��I�^&�6J��ή��Y��L������i%i�����AX���8o
����`h�ZE0�+wT���a^�뫿�~a��J���Rﳡn��_ݨ%� HJG���t�s�l��#sM��A�u�0)K�X��6��´�aw��'�)����s�s_s� ��~:�M�4+V��?�������-��Ϣ.#;��d���(�к�Z� ��wqL�}e/o��/!ǡ����~/%���H��a+��o
�Do�-B�k�$�y�_���C?"��o&��ڔ/���_���Po��b�6�� ��};!S�ũϹ̫�hk&h�~��PZ��#��"+D�&x&� � HQ��3-r`ޫX���W�$��yƉ�&��d�p�u��IH��Rϗ�h	F�\���s4�J�}��'03��@1d����|���|ݬhv��#8'��
��(�}���P(9*�>P��`\�z&� �w}e�:3.��X��5�K�X�{*�C�{�x�N�W-FMF��o.{��V���L�N�U�XoJ��U+�qG�ndx\JK�V����H�ܿ��6� ~ ����t���3~�;�B���J]^S���55�5%�޹��*l��U�"��^��z�Z�tא�CݨEՆ�F��8Y]\�pk>��~�����F�9Oe]����ɹL0�x�ܧ�U(@�@�.g�]�-X�@
�:P�E�����?sq�m{E{f~Gm�_���3/�:8�k4�S�N�_{��ZJ��z@	��TX�-��h�\r�7e(`c,![�������H�78�Aί�p��{:�s�>�5���0$����w��}'�Ԥu�\!_M�j5&��!� ϱ7R�s����0��ot����]�֣�\��p"��� �'�D�Ng>Qԧ'�~l�6�B���﵂龜mA��h��k�2�Ǚ��jQ����a<s�Ũ��&�H���������W����3�ȍ�E������[	y�)���~t��s�l��l�]-,xSQp�ި~9; �++�m۫p�G ���y�m�#�Q�HHP�i�d	Q(�n(�EЏ�OD6$F�E����~���R�s�I���J�z̀���ڐ��1R��lK.�{F.���Ԕ���6鲊�?GZ6fƧ4[їU�_*%o��4��U�H^ڥ�z5�MC��}�;1���ŚM��:!��ͩF�yK�c�d��-��R_U0����2~�Q@k�#<��}�fSMUHxs�1=Dx�e_r��lQ���K�ƢBBl��ф�)�$���,��/�J�FW�^6������W���`[`�&u=W�\6�&�Qpx*�Ulr25Y��I@��I�������t6G踒K��h�yqP�j�]�	�]�3��.z��+^���J��{�Ho�?]̃�b�+v�\V"Mݜ��ѴT�N�lv�� �dx��YaL�M~8�Jw~��G�̍VL���r*�M��r�6�,��d��M5�q�L�M�c��3��@9[b4рz!Ea�-���W��}`���Qf����Ⱥ��x�?���E~��u���˸���c���C6��Ja��^�	�J��۞�?|�w������9����&�N�[PEJ��7P�0���Y�[���o��d���0����g(+�h���_΍��(�dA�F��7�}C�n�GY�9dEəEr(�s���r���6Vr�K}�mF��wg��kL2�<B���Go�
�J�̕��وn���Vq0�r�ne-�Kz_��m�g��愝|u�KF��kAV�m�\��YV�B*܎re5˶�%߳�V�4J��Q��Τ�+9���6K��Y�͒��o��L�m���y�M�MY��AnE�D�k��w<�k�-Ϛ��n�V�׮�NvK�jx�Je�$���W0��}탵ɡ+D�;~��v��,~���Gv�A�S�(�	�iw��G�U����
�z�`�!�g����1(^Y�\�u�a*���]dV��p�=[x0/�W�RY�gnL�<��^�M��)�ӛ7i��V}.�!�a5���}�lS�;��)} -]R��~Gyˋ|��R� �y~�p�}}3,zʘ��t��r��DE�
r�ס�9�P��m�䇅G�zj`+9Td�?�Å�غ�5�6���ԕy��f�viPS�4�}�`��E��R�Ej��<��\�e��l���)�J�}���R�`��K� ^������jecl�8�2'	|�B�)��s� �n6�h��~*��콚zl��G�X-#�������������,��C�;�ġ=���'1dMqna���Y��3�s�t�O���w^��x�����Y�<#v,�%��s��WL��J�j�z��j׆/�Sfр)<
�7@N�������ZHҞߎ}fv��NRv#*�F I�0M�g�J���\E���2��Eg�2������sOȇ�+H�ý���S]�؝����6��Q-h�N�BҌ�������I�M0~�a�s��^2Z�(�W��t���J�m�r���fQnj~v�׸�ӵb^���TOSQ��Dt� ����m)In��t��s,p:{jO���l�5���̳�L�޴]�ö�M�v�>(��K�z"
�U��{Q|���e��H�����_�����d�?�d�e)�ܢ��)ɣ��b���]snv���h<���4fR���uj�����8}7I�g��*i"D�H��?�ɕ)���3=���lh�e;Cu��4m�H�r<����ƀ��#��S��'��T���C�mc�|Co�3n�$�sw��.��k#��x<.��h��e�φ�^���+w�õ,����cW��5mJ�i��Jxݓ�ya��w~om�jl��|q�CG>fn�I��t������K׏�%��*�M��X$ұe��G��oW�3����Ty<����~�5J���q���1�?i�T�AUE!tJ�k�ude���$.��;����q3����vQ^ �'E��Ez��&��N�&�rm!m����5v V��	�)��5Ɠ����?Q#�;�^�x,�<$���E�e��a3G4p��<꣋~4�
�z�k�sf:y��YL�ԈCg�d���#0��My�i��t��F���k�Q�N��"�tc��N�+�P�i�w�@EѽU�c����W�N�J��zg�%�&�{�'�� ^ަ��-��Eŝ��-�KTU����6s�G#mx��2 ai���Q7��[{#T�G�KtYt���iojx�N���y�?(O}�w���/�1�1�I��W�ѯ�Z�i������,Ĳ7
�W��>��߈�|��LR�����>�
]��c��ΩZ�HSR����BwS?�O��S�ّ��!,pт']�x�!,�#�D����}+i~Y��Βq�N�&P��Q�׎��� u�ٗ�)��?�~����@/�(M�/�u�v�Tv�?T�<BW�"�c�7s��1���(��G�y������o�+Kr�/>��KwG��(}� h�X��H_z������T$��7�X^�xޥڮOw5�t�����,]�T1ѡ����-�-TY�� ~h�,��Ѥـ�,�A\n�1�2�~@�*��%�P�Ł���\�pzij�7����Mu���u�<�pf�f�v.���
q:
:/Q�ȁH�E����s�e
H���8����3M} �L2uk�6ߍ��H��H)n7p��f�w�����.Nii�ﲙ{���g�8���%��3K5�x��Cm�K/]Q��@��J�:��!z�ӄ��G�(NS����^u��0� i��@�SZ��R/�s�
���7��|���h���M�߰�
�ǟ�^&u����N�@�0=��ӷ�;lǙ��PM���_ʩ�]���Q�!QQj���v*��Q@�eTqD��8l�*g������h��l@���x���5zᡧU8I�%G��:�w�GLN�ݖ)��T�E�Rj_��|���c�3O��MNǟ+��~��|0�@����D�0D#�)K���V���fX�S0L��Vv��KU�e"�/vQ�8w��KV�Έ��&�L�?�Gb���3-��]�Q�g;�KL��q�(�(�i����ڞ�������Y��29����û��A �������Ϭ��7A�&u�oѼ�GLa����������ߑyձ�A�y�)릏�8ʒO�J�Q�Ǝ�] �����թ!B���}M�]��^ZI:�=@O�3�)/g��M�����`4,Y��lӨt�nBc�����C�����?���0�s�}r/aS�� \��	j����Lw()
�߬��e�ţ�
�N���\����d_����wg���pI���(S<"�9�{R����X6�WR��	˼hO�sh1��4�G�U��M���3D��98vZ�r���<u��2N�HWx��"i���4�y�c
�_qَN���������;���T�z�F��q�(f���d������Oe��	�L_��/�Vy�w�vH�歯o�^�s��֦�å#ػ4y�I*���ӾT)|S��cK7�e�R�ڎ��9����O��\�b��&7���E�Y|���w f��z<�tn�0���AN�hǠ�� �=U�MRfɧ�EEMA*��rIz�å�ٵ�T_�*PU�T�m��zk;(��+��.[�A���e��O-����U�ӳ'�O�������j�pݕ����*�u�m��lC<mB�A��xe�$�C�aMܸ�3��U�ܟ�)�>�so���?�'X�V�+��Z%qM���s��lu����0Ov�����
���y6/g2�o�U�hqE��s�¢I��� �:���Ն4�R&�\O�N��3�yD>�jV-g��6L�|����5$���(3������~H�]�L\�\����w������LIIab_���s�_M�_��ܗ���������A�DW���OiEΜ��'��u���hq(Z����{�������Wqs�[]��g��_H�x��:j{�Ez�5!�6��Rԯ�<ˠwu�֥��h5iL�h��gJ�^k�U�O�oH�P�4!SE��)��w�>�n�� ��#^���@,O[�?G�'>��P�-�1ku��6��&lB�%�E!LJ�����Pa�Q�?�?��:�-���7<�7�R��f�E��d��.�}~Mj���U�P{=;Z3� {$�ͤ�܁���X-7��Wm(��0ZS�r6�n�CkȪ�2R?S�f�4?O� ��_$�����a��3�zz�㐇'L�8���EБ	�`�e3�� J��+W�����6M�ڳ�����k�N��|��Fs�^D����"��C".��q��Ϟ�q�ʞ9������\��=�E	�g[�
�����]_�V$��eѿ}i!��:7K��Xj$��qB�R�:�[����O��فKUß1�Sm����MYp�J��p�l j�����܊�É�Mz�X�Զ5�~��D�e g_�u�������N��P'����k8`���?��z����?sAd����B}�xl�.{KD��^�\��"%ʒ3�|%�YӠ���bKJ93$��OV� ������nkɿ�r��fy4�N���R�~����pIW���c&�7�
�곡�<|3ca~�PM�
�nz��(Aw�G�ߪZh	A	#�f_��B	�xh�W��r�a�������^�r�/�Lyp����&��?F�迿�Yݮ%�Z ��Nqm�tQ�#���'�~g��Dֲ���uS���ك?V~�  �?�3��U������/�w���������9i�G<��z�ո�y̓�~��c�#�^��_���i�-� �"�8�<Z����ܾ�����2���v�)�}��=�#7s���ȸ���Ť�il?l���]�� �r�wa��7}xo���* *.��s�N)���v��W�p��$�����/�r������M��NK���ߙ�JW����Ɨ֖S��ca�r���Nq*	 �K�
��e��
N0����Q��6�&$�.� C����k������O�·���Rƹ��K�����)QՖwէS<�K�k�ʛR
�v�J���9r�!��E��V��I�|�@"�ن�1�wBz�.xhG��dZ���cW�e rO7Q<�x_�F��I��Ley��@0(⦚�˗A���Z����ڏ�?|:f!�����G���'l.���9a(1�G��x�J�q��L��5�!�P� �ͲNH���ف��1�?}�񡱿	k����6*ª�)��o�S d�LL����fi}���]�K�@��4>����B\��M���(��y�D�gmB@��<�2̡[��U��*��`���ǳ�xo���o��FZTF�;N�����6O��e;;���� ��5VdI�s�r�Q) �	������T$Rk�߾�cC���0��"_�g!rA�;��A"�o6W��=�#Cc��JR���ykW��B�/��G���R:��w||�W��U�˷�E�'7;�/D����rz��`�߄�C��vf�b��ݥ�&ߩg�J�B��v��]�L�&�1bv`��/jք<�4}��pqc��T�)I�l������^u�$�r��ed�`�,����:vzW�I�Н>�W/_%6�"Щ+�ا�v�1�;oW����e
����A�RC�x�d���v@g=�j{��=v:`}�Az[ڗO�~i������3 �m�nH����W��Eq6N.s��,����-�iƋ�+��~�D�!��F�c��>��@AN���$��66��UT�8���ͬN�'���Ҏ� �(�vִ��.���? ���|p��/��a�ۦ��YY`2)���/�	5ɝ� f�������ӿ�����"�mZ�
�ޏ�.eK@IE��d�ľ��rY��^�i����]=���^c������ǰ
.�v���F.��p#�����gt������9��7l�NO�[��e~؅nHm�13��)�@��M=�S��m}������$U��R�Y��b@Oj�ڙ����~�;��q� �u~68�������i�o����oܻ������ܛ.@�ӌo
�\[Q�Q�JXٛ�^й�%�G�l
N1a׮C6v8�i����y�|�������E���E�|�F�EF/��7�<��ow�Q���t��!g�"�o㲿P��4�>t��u 5L|\��!�m�*v�	�O� I���Y+A��+Qr���e;+q��k��Mk��$(��o(d2�� �A�f�ٮQ�g�
]t~���b�§�]0���WE�߱�Q�<A�E����.� �Nvq���` |��������##����@�A�6%1 t �������'w���	� �@�VD���y�R=�H���K�=&�;�^�n�.�S_��%���{�y3�+ʘ|T�#���-0na}���~�-@wF�	�L|� ��M���2l���:5�]�W�e��K��}�C��Cru`$���z:������~
�=/�)��r2��2��x�h�t�;� ���x��5�*��\�Ose�$���Ǟ�� �<�sbqG�	F�ɕ,~��\N:�w�3�	�;���;���|x����/��o^*��f��V��N�Ƙ���	 ��	{J�j�SH��Oȧ�m�{����Z�c�xJ��O�_Ew��쫡�Ɔc�/^�}�����ӵߛ�Uq�:C.3�����A�\�ځ����*q�lU����$죈�������L�>�Ǹ�`˾�2�R�De�-k��8wz�8ƀ�V�l*�͏ ;�Pv��I���}�rSX�KoW��P���Kc��[�n��@S��}��'��`T��Ӯ�X�2XY���ad�{��F�� n����K^"~�b��j�/rۼ��\&4n,J��؍{{.]+{Љ ��o랴���%ȺG��F@+(WY�ӯ%�Ł>�ޞe�э�_e0��C$�C����7��F��~���1d��K�͖�Q�� �!zE�蜝���|�����6b];�]W4����?Gd�� t�-FE�	t��U�r�B���d����l]F�Sb��j���Xp���,+:�!IC.Ȁq�L��~��S��8`j��~� ]WnO&�B#�>��sY:�N>��� �((�н���F\St���EC{kk��	��I�{5��h�Zֳ=:��()��$��ܒc�>������	���'�["�PDc�>H/�����B0G���c{ɜ|��~�c ��4�)ū>M$&?�����/4����2t6�e��>���|���B�e��rf�=wZ�����\��h�b5{�Όww}:��*A�l��`�X�|�j-ɢ�x�nƥ�~��܎����pEA��IF��}{0�� \6�8��A�H*KU�t�`f���E|!;�^F\���/U����Yϛ�:Ƶ&GA���I�TT�΂G�99}>���>�q���k����;k������B�O(t�l}y<������n��n��H�,���5(��}m����WeʖK�*;YʾO�f'������Gx��}<���3����y�g�xfn�*�-i����O�d��d�9t�ŭvB���S7��L�\������m�%˶�*�[�r�̶�JW.p'ik��7���b��������Su�
������G�K� ������ь�ڬ�O�pg/n"]�)X,vj쨍�C��V��8�{x��N��o��>|�a�$�����8tY8R\�W0o$��r��cp�&Msl��_Vh�=�rT�z����2{Ƌ�p��+Z�!��+��RS@�����6�A��7ݐD$�b#����4ǚIn��_�������ۘ�vW�\N����KE��[u�iƏwH���k_M�l�h�a�k�]���TnG��f��+�؎���"뜶�Q�U�����ü t#K��?tˆ|.Qm�[8��s ��+C��VkvUnb�$w��Y��=UA$�[GۀP?��J�
TDٽ����KJ���'�NU괧��iQ����@-p�����I���4#~޳Y>��|e/?��=�aoI�s�.�a?�苾�N-�w���t�;6��s*�����0�W:6d�J��{�:��h|��'�)o�s�H��k��\�|�&�V<�l��/B]y?�Tae���8���0�.��#��؆�O;,NB�������B�;�?�gO�a��N?�n;��`\go���ʒm��s3�5�.K�f���u��m�����lz��5��"��Y7t���p��ħ�Kb�e�Gm(��/}��"�芍t���e����o�~��d�CP �+�8�n,K80j���n�o�tz��T4�����̹l2�+�➞�|�{�g�&)�q���a��v�d�a���D/ǿ��G
�f̷�I�f����ݪ��Py���������w��|����:������:�rfT�����?|,u������쩺?I���@0Z4���"
�iQ� �tC�i[���Z�1x�� M�捙L>݀�t`�^�lL���*$
�.
�W-�6��Yoa֙Y��EZ%[Xr=�̣�;l���΍�X�b
ȃ;�-	�_�oԎ�?��]�Bq :�����6l��̥�I^ݦ�K�J-%D��m4PB7�[��O����x�>0>s�ze�L�F]��&�$�䓀O6egd�ob!��*� E��b�7	}3�����P(��(e���NC��Ҫ\ƨ���ͭ"�.�¨` ��᠊*���LAy��?-EK$��YC��R�m����^�v�
,�y�$؜�P \RUxUȧ6��b�5�rk�ĸ�B�����;�j�=2[�c+�j��J�a9���D�5��P�}������MA�_BF� y���
i��	�&P�P�pڵi�%t��nhftg=j?݇I��H�� ����ݚгqG䵝ə0F3��մ7
6#W��@~p2_1�EY�6[�1���֮.yn�m��Գ,�����_"������4���e����,o+m��ϥ��kf�71�mL߷��ߛϪb�`!Ty�U_������j�w��n��u��d+yZ�H��	Wu}5}��E���;����X�_�y�j��J��~<�@�?����_��Ɇ��['M�Ic�C��0o��Z�<���f����w/@$I�������o�إ����E��̆D�f�R����;DME^���l���P_Y�?��W��P}��ۺd�Do��x`q;!n����ڄ�KC�o��q�~��)�6�W�pi�� �k�	�(�P��Udppr��U����Fw��:�k�/l�XX���M���_���n�Y�����v �v���a��;��y�-�`ڍȬ��*��[������5N�C|{��A���߸*�n!9Ԍ��`�;�6{}�!ea���ŏ<�8L���U���@��뇫Ng����j]��Q�q3��B� �77�0��#��V.e�@���Ϫ�[xD��'vG�����4;?{N�=���(�e�H�r����G����UzE����me�/��������ќhrǙD,�V(�m[�f
[��o��r�Դ�O0����C�(����6ow��@�yU�:Q�*�)�(;7�ޫ>��31<3#�b$m�3T��)K�����c>�����$���8k���9]�6��mx�;�����#�UT�l��{2J���<�+�ױ�W�/�6��M���|D���(Eo�
��1x-��]�E��K5/�wR�q%E��$��ӆ")C��贴�K+i:q�"�i\��&O�����m�+��/)J���'��+X�Eҿx��k�Fڔ�`����c ��2�R��t4����������$�a�@h�RQ7���Q��۟�y$g�OkK8ľU<_��ZX �0Lp����[R[���ړR3�&�C�'��U�eo�2�:�]��=>���B묬�,�1���Zl��ui��~�6Ȑvg�ٌ��,�"C�C���������
������_I��3�(�K�f O�	�&���W�AŃ؇�6���q���g&�����2��辰�[CB��r�IwxA"|w�֟sfd�Y��v�����aS�3gzk����x������
����F>��/`W&�b������{�Z���p�ܚ�i9ޕ#_��Tg���I �u���܏x6�ȣ,��Bb�3wވ;p <WCS�H~b����݌xR�rj�C���4��]�bM0d_Z�Zfgwr��xǖ-s���£���]@[�ob�'+�;tl�8w$�Z�͎�8�o6����!�z� �+��� ;Y� �A3�Z����q�!���v����ғ�"o�I��Ԋl�_7nؕ��s���	�Kٍ"�*\R]�E�S=̩�;�O�&�V.��b���\|��U���t��g�ݕ��D3^��9�FK�`9�Hڕ���h�L�P�ڷ_<vf�w�9�ʜ�Mqv�F��k������T�Nt1��;<�Pi�����I�Tx����
'�!�M6_���Lq����\sw�*�U�f�'�N���{�Ivk5Jo-|�]�F5��+\ý��T������-7�m�n2`e�(SX�E(8��?ޑ�bN��c���ħ�)f�~�����4Yd�.��~���-󔊷|-��K�*}(���ii�*R�nK�̎Ō�������jt)u]��.;V��0r�*Բ��U�9��t�io����2����v@4���S�M>g���4=�˴�j
���霦A�j/a�A�	y'���	�����	�B�r�5~J%�J���A�j�#�%�yR=`���j�Z��j�Iu/fi%��z�͉(��0A��N(��ve���'�#. =��sٺF�C#\L�}V�a6�xp���i��=ɱ �i���X��&`�lOt��^Xt�m��Y���8�����o?�n�<=(dm�@<���`e�Ӛ�gZ7���	}�ϟs���&�ff���/|N��G�Y�0�5�|q>�ȱ������V��dH7Ӡ8ˤ��-���E� �E%�{'����t���W��g"S�=i|��O�<&��O���ə��_���AD]V�R�����,����Yd���?��ؗ~ �P^+�A��?- �-���7���mM�HS1�@��y^;0�ce������޽4�!!�-��gẰҍ�N�};;B�}	��Q\*�g���W����'��W�a;sx�2�-�P}׍��RNK����C8LS���ꜙb���!��J�� �e��2t2WS�����旁�bsCv�[Z��ȥ�X���ٟ���n�H|!�x�*_�
�]Ö�q�_P�(i�������$,�<"�~/!K��բ�_�_����C�}�\�ۺ9��wT�M�5�����@�W�N��B���=e;p�<�S�0z�,�o�5����bQ�v�|�s�]A�?��U�-�2)��\iѫh�\��N��z�UA벅������瓴M� C���g@?X?ه��~
N�.V��fy�k8���'T8˳���0w�*{�u,~gC�C��w�9s�G
d�
�g�T�d�g9��DG����ò�C���\?�Q=hь��c����0w����Y��z�a�kh<]턾�N�; 6���[��ނt�f0����(����󌤇v1�03[&�]���E��9���Ho҆\���h���V�f˕�����x7)�)��y��u$��ts�Ɨ��FQ�v�6�ً�\o='�̼�/�l��Z
>]ݧn]8|W]b��J&���)�kwp���sK6�6���V�R:Ս�cdT�'����D��6�9Oy`�� �]���%�����Y��N�W�h��ogh�9		���2��Nn�R��O�fQ������kz�Ef"ŷ��Rh�U��K *�d���М�X��#�����j.���7J.�	�k:Z�O'��?h/T'�����S��>.8�8AZYF��,��T@�N猙����h��G���OLd�Ep��N]�A�ҕ��z`KX�;՝2�K�nR�pNhK�E�>��4�	�۸�Ӽ��_9���ci?vO�j׉��z����u� c?�HP%�f�{_�&�!\����̽���9��^Z��O欧9��Q2Ni���W:�9o�OT���s�����wꝫψP�<�M�`�*`�|c�@�n���be6h��9xVV�L\;��r&�n�B�ŅN���g�@��5X�n@��ST��&$���>.��9||^�S�6,�"�[y|5{�s�gƝ��q�Wq4�ͦ��0��T�,�?յ{_־U�)�[*4�����v�e\�H�5Q���߶#&75YCF� K�J�bG)ׁh��Z�,�i:��u
�\
C�*%xP"����iۯ���>��#a���pw�����7y܎XM�h}����=?���uѷ�/�@����5�w� �Շ��dq���~��6?�̛eǽ�g_7ˏ�ׯ���8�^Y�B"S���8^y�4�� +q
�L�X䑜�s)0L�G$W)5���3w< pn��:����gq�-ݳ}䪾�51mr�>�Wc��!��1mS$��`=��������(�V
f&'�k'0ѢT�sj|��|}�"���?�B�v�/[�=	{������6�h���b'wIY��wnI�f�#IX`��i��`���O�X~�ܵ��lF�,��-�3A����8%~����F�~��������I7��`���+�m�j��#�R �t��:��V��Kf��L��3��A�9���Iv�r�_݀�*k�j:���"�J�5�����j#v�F%Kp����؈��Vڽ�Cê��IW�Y��q;P��7���>H�'I�A�~[V
���84��-%i�MTbpL������~��mu�MS�մ�������Gj���8��/l�GZ��S1�g�_Z�4�0�LC�'�o@]¾J��
x�w<�os��!'��?��斖$����NؤFn��ɭ�p�V�@���'nD�oЧ{ߏ�07/8	[��M��0�X�����f���	Yr�h a>l��F8�*.�mw&���-hcC�������;�X��T��pd
����<��\È?�-yݝSg�N��=�`D+����"y�{����ok��7��W��t��m�c���I�|ŷ8��i�R��&**{����I��_yf�6�r��:�ف3�ގ�Q����3i�i0Z�1�L[7�� ��D�;gT"�W
�)���'�}�@A���7n��Gv�1��B�
�F���N���b���_�B�NG5L�C�p娾�5%u����O_��
�����QO-O� �9�����/�^�mf�'����M�M���3��Cg�\d��OX�9��Í��#�����V6�tU�j�����9�T��V3|(�Ǡ�q��Hwg7q&ŧ��D����Q;�+pSgSc��f�}}�⁢�ax4P�,��P�C(��'>�C8�T�$�k��	�F~��@9�4/(��A��8w����7n;�ZB�����z�v�!��Iz�t�Lr?���$H�A�/�|�2��s�F|�Z��Sz��4`Dc�������'��i^_mj��Xs8�/�m�-Q��drZ�XC�9>#5"g-Hq������W(9p�W���z�4����P�9�
n���x���T�%1ZC!�Ձ�/yӗ0�O8�n�}>����1B�ڦ�|�� ���Ž��{�iG�c4��|��FAW���|<�ǹ_u���C����45�Oݗ��LM��}8�A���rQ���0������"\Nr!�k���k�绛��M�*�c��X��䗞�+"�zfeqf2_���bnN�\�tOgh�pM�������J�HB᪷�z���0��9x���`:�k�~݋y�����+k���sx����n�ب�֤�;��$$�oi�vWD)��6/�j�
�Ҹ'�R��!g�"�A	uk;�i[�#*א<�9q�)�L�>��DCx�֨��b�{/��e��dN��s0�UB��6�>���Z���OQ�m���>3%'��u��H�%
p���r�m�oi5�˾�A�0���;M��)�����sh��mN�2��?��ćиó6��נ���<��-� \���[����|P�@�޸w�?e�7d�(pղ������p+��;a\�P����y�����㲻�� ��0�� �m?��+�g�)�V���a����V�f8tr�s�����:�Wt��gՁ�}A���2#��+?��{��ni��cQk"݂�(Tv @���16`����`�.���y�qvl|,�ߤ�rŌ9�U��:��|��/����`|4��a�I{��V0=�x.�J_�c��.�Y�+��A��i ��1���v@�xTbG�m��Q�7�v��z��8���F�Yl�b1`��t�}�AX�Wb%Լ�C0���[ڥXjb"_�{3���R�����ZX"=X��K�s5��PP@�0ҋ���
_�s��W(��f�ὴ�X�q>O�~�!g�0m�swSn�}vAf�l��} ��z����%���Q��;i&Qv�߿�H���A�G}|�Z����_���<��\�>��:
�Z:�)̲�0B�t�N�V���.ˎ��z�ͯc5���l%m�,�&��3E`��,7���Cx:��Iǘp /_π���F�/G�]��WRv]�k�[Zvd���d���g�,G\�`�c+��P���m�5&Q&穳ީ<}�]xX�>�tW�,��j]�!D��_}L�R`��殂��%��f�����kï��$�ēL4�y{�-�.�'���?�+}�;6-hU���q��ب'��Xl%��D\8L����vj�9�+�*R�X�w@ t������ؤ��չ��JeZ��
�\rf/Zx0�:�{�w�<c��PREǉ�{4ܷ��N��g����|�j l)���Pc��L��f����\2��q�L�WK�����Pg�9
x�����BJ�n�6簗 ��xU%([G�`�Ţz���6�&�g"�nv��I��<]��_O�J�-S�QfY�l�/�
K\;�%H:��U+�QD�͈n�>��t�ll��f\U�};P�Z�W+�,��8�4�nT��As/�ݾ�O�g{ǁgv,n�g�u�����	Tp��������R:*�<.]�,Wy��b�f�o7�?����9��iu�b��W�otQ�.���e�>�(���4������k��F�m�-��Kx��Y��9���vBUrOiN��VZ��x��������S!c���8�_�M��#�}Dx̯t[V.H�����Y�n�]q�����M�k��H���Z��������d;%9P-�((�ܾ;|����\q�>���,�ȫ���>-}4 �,r~:�
K���$�f����80mѶXv_nH�nv6$���x����.�+q�j��j�J��A;���Y�	
����`�`Sf>��ǆb�Kۤ�6o39�kɦ	X��)*ui.�/�o5���b�b��C�jь�<����/�K�?�+�ރ%���=�B5�9�T��4㐴7[hK���8k6Po׊�� wٱ��1ut�.�S0���Rz�3^Ld��1�q���#v�-�7/�����g��e.v�U3�R�;`��"�-��cu�ͮ��WT�$����Lw�6������]�YZI�����i�z�݊)v���Y-W	�o�����$:Ty�b�;4Y�~}� Ň� ���9��~�ߡ��Jͱq*6�h�̞���>���1�����$ԓ+4�|��h��\����2���C�è�>�MП5�ּ�D�QÂȔ��2gA��Ǡ�^���g��"�q�]_��j�%@��3�����O%@��J��Z�W�t���@���F�~{�U��'،컡@u���UY���0����"}�z���v�-v��&�x-z>��(?�����ˊid7����c�e�,��)�L�,�������Lj��U��#l)�UIX�n�H��	p���#���p]��*RP�u-���'���(����QCE������	>����!�w�.=��im�����Uq���ń_�v��2��w�7�#[%��G�5�P'n9� z��F0�=-�p�����a�f4z���\��\�q>Z�d��sJ���D�2�,���+��)�F��{VBGM�,'P�� F�8K!�ޡ���3i����d�+hA5�U��F�s'�,�l�����y����\?h�IB@-x���8�[��\�?;D��HnH�ҜoܧZ�N���B�R��:�E����4`P�����{�Ê.ptdp��v��o����'43��a�*9;t�r$-���ޥ{����y}��=Q�V�D��{]�u�w���3�T�r��@���ipX�}�����
[�6�.��YQ�S�S��H��f=��kϽC3;:-�t����]��:CI�55�N��pw�A����o��'a�;u�����ǝ!��w8�#1��#W�&-���0�B��܃�:C_U�r�~p�~Y�Ǌ�6TU q��+u���\�/�$�j�sBW���Q�Tj�}#�b>����\@�T�X}g��on�"-�&t���~����� �
@[;w�ӷ�'{�"%-a��������*p�u��I`�|�P��ޞ�U�l>HT
��F���������ˎ�͇&z��V0;�G���19~o��jB�;�a3F�!@��h�p�TTû��|�6����	���W�O�J,;p �Ȥ�������iP?���.�y`'G���:���m��_���wf�-\��t�Dd������Jߒ>�(7���`m�d;x�Ր\��ww�kQs��9�B<*�oڧ�/ -�Ai��N����z�s�m>��$k���?��=��N�� u׶�<���s���g��ڟ*Jӎ"��@s�`���6�YU��2B>9�W��������eg�A�h�d��v����l���>`�ׯ[��+	T�z^��~���d�5.��^�3^��V`{0Y�x3�jXw�I:(�^B̥q uo��4l�E�����$f_!$��?(z�t��|���A~���C az�^[#NʳMz>�v�<�܃���\����o�&/��{�Δ�q� 
]{B���#a"�|7���\W�Z���E��	A �<b������P��M��
|ba�P����ǖ�60��w���̤�ױ��F} ����f<b��
&����#S&@*�h:�	����6ý�6�1�*#���v�$���\��Rҏ�<T͊�MQN4�e:�e�A�B� �����FA���!:�3��CCcAOq8��4�geDu��\��E;e��c��	p�����Vo;�T�KDЇ�n�]y�Q��|��j4����#̭�tª"�SQ�a���w��zq0^ǘD)va�`���P�k���9�^ܘ�Fa�N�/��N���p�:S�q�
�1�pvw��e
��0N\��J�7l��v�\k�MfƲn7�4 Ǯ�͈�b�n��6�g�uX�7��鯒'��o>>�n� R[���
C��ם��y]����x��Y����u����E��g�f��+�c� ��_���/d�T�Z�J֜�6���;�;�;ave��7�+�@��Y�~��� �m�)2qUK ���=��:�+�İ-�8p�uLH7/��y�Шo�H��$N��dK'*'���#��y��{hWPw!~�
�c�`��#S\��+j�QN;-���H���1Em�
��3Ǟ�r[�V~u�̽_�vxG�\�3P������⍝TT���V*lʦ�G�a�o�9(��:�*:��
B�;��Gq��<�Sț]~���i��*���s�*q�j�[u��D�8�v������$�n�S�*�Ӻ=٣��ȧ��^}��
�q¸/��H����p�_KkO�*)Q@��1�&�L�W{����x1�J���\���	8T���~���L�0�N+ḇ��z勴G�mXPj�Z�<�(v���*GB�p��ud�����H������������x�A���0�iO{
ļ,.�D��|���@�J��R�/���N�i�Nf�Ò��hgnk���a�*�-�!�.�wd9i/T�e�@oA\8d�ċ�������H��.�]�UI�Σj��8�6E�1ĕ�ۊF�#K���U��a[͝���"oow��5.�Dg���4�>�W�t��sƖnD�\^.YD�[�F�!���^	Q���n�cs���$�GÄ�9=�+��|��$���7�gȴ�l�m]ֻ($�T×�w:�����}D�2�_���`�V:NN�/��F�2{ˌ�e��5���4�15��o�)}1��qtI!K�ݐ�;9�F:\c�@����|�1b܍����Q{��:y�}0B��X\Q�!�s��By8�,J�����%i��g�aR=Uj PrKQ��srt�e�r��H���p62�'^�,�q��N�Ve�EStz}�ACZ�k=g������K�����u�]��w7~V�;��و�o�N�"�k�ŭ�����ŜR��/h�ן�t{i�5������<a���ow�W�j\��{�����{�ޏ�g���"���".�.��A_�b�x��'"c�����G�lQT_i�u[�k:�Ql.�i���־}�JL�������FA�d��Gt�B�y95��l�p�ڪc��l�?��;�ޕ"��_]L�6��V-qw��%4������>�79Zo�����o�T��	u9��FQ���>�yi=$�ӠT�ɻ�q'����ҍ�T��!{'6E��U�ዾ�_���M��Җ9��U-�~���ǳ��j�(�1���������j�\�9�[�D�vh�)�o�G�bg�E:�I���uF�h3��j�	�o��%���@�:6ZĔD�f�궡�S�_Õ�ܦ�8�۞���z����"43��e�^@\'�b#������o0З[/t`�8�U ����z��ߴ��A��l~M]�1�>*RaK������ƇG�rw��A~=�8wa�+J�S�2%a+�*̓�'�L:P���n�A�2�(����G5Eik�� ҭ�&�Y������yl�b�U*]HlYJgqX��XW�<�%�)��Os�*)��z�Y�V�|���z�K�F��LB�r0b]�%��/�~`��+�NƇ��+���U%9>�ư�4�Ң�8�Y�=��]"@�X�Y����N�_�/��ԝ����~F*��6;�qpАȰ�D��z}�������������P�E�n^��
~�ӏ$�A���$�?{��֌xL����cל���جSRq9\���8�Jd֐�H
u5�q���N��G��Լ�8'D<�fA�=�b<ͱ��a�^�}��jb������Z��.M9B�c>��_�F2_�uM��'fQy+���.,m��6�ġ���Y��<����rTm���XU\6ΰ�*���1�g��<%%�kv�4���������~���k}���e��%�����/�t�5���O��π�|�_�>W�VEpq��9���F\��UO�&<`��B�Ȅ�Ԙb���_�tt?���O�!�Ƙ�9�N���a[&7�_�Wj;�9���k�h�0U�̾�j��f��&޿��8�Oc2���*���1p������O�{�b��w23��R�������U��K��l��G��Γ���Ջ�(<}2G��pj/^��SAh��U+������d+0���!z�u�o,T�z��r�;����L��᜖c�o ֔.�^��]|�>s��̬��⭝l�;Nւ���^�o��e+�!l(�x��11��L�'$�nj�׸2zV�F�����ꮝ׀��A�b�fo6_F�d#��U��wie5Ե)=�7��AW�.7譔��D!�`��CcW���B�&����|}0���X��Eɐ�H5��Z�48���W�H@D��[s�;{K�T�k&:HX%�
^����=c���N#,� `, �}�gb�tԔ�O�m�z ,8<����Cf6�)A~;l��F����6�2�͏��q/�x`���^e�j��a�%o�~h�TyVJj?��6zN�2��S5�!ș��m�w����=��	T�q>oUo�����W�OG�8�����xi�d��gIgR�S������ٿ��ԊZ���ls���x?d��Js��v��j��z�Q���ո��>���n��@I!䃹��/-h�|s��BB�U�;��~��9h^�b�w5�p�w���NG�RX��1`��EeǇ��DD���kP	��}K��Ց8N���ͥ�+�a�����kp�4�0u�[�=o�'�����98�a����\��C�}���4 �z$J Z;j�������������Yo��H8}����5��c�k��������9QI������K�"�s�<sA�E�x�X�>��"[�v4��t+My=�����\/&�GL'�f�����{�`����N6Tg�|A��B#���:c�)@Y`��� xYŬ��D$��(���jk�j���¤�l#}�ʠ���D�|O��^�c�( �����a�d��KR�Q&H��9�������{���u�E��Ѿ�V��.B[���f&���5���_�U��S}�4�D�T�ߋ�_;Z�W'�s���C�rz�?����
= ��J@�e�w2Q]=���'Rs�u+8I�Ѩk��*	�D
�T5qfT1�(���|��Ϸr�ěO V�S�$����ːf&xr��;h|�i��q����I�utt�iF���Z�5O�XQ����� �	#� �I<5(r���@��'��h](�}yV��֜v��[�������^m#�1�b�x�?}a�E'�5�q�-@�Dob>��
̷�7e�F�F����ݜ!Ȧ	��O��p�DP�1���:��~�:�]Za�ʹ��J�v�KF+��d:��D�����eiK�E?��?T3�`$H��՝���"�P�jY��h����8�����)kk�g�V�u�e�_*��3����޼���=i)m���a�-442�Lb=��Hŝ�}��+ (����H��H�������sz��S�p�C9��DDXg5��m���n�Y��QK��%�����jͿAj��B�{_>fo�N�T��ֆ����գ��8�S۟���5���&�^���d �V
=J��n�/qUg#���uk����Y�夐O���ȥzN�\]��(����_c�@+xP�V��ޫv8w�7���?�땇�d䯙�h���%���uiQ}�
5�?�7u(e����;ź]��L����1�w�B�;y'�~p����8�'��l �j�)������4vl?�	X((,m�Z����^�_~��*e��a0��+ P�������H����̚}G|�`@���GN�t-�/T�N4�g"
;�L��z�����	� P�-�H���}B��-�\�_Sc`>����h饹*�A3����9&��i������A�y[&0��a�
(�'S;��ّ�g �f �8���p0���	 5�T5D%��c�� �.A�J��e'�Sl��*��P��D��R��wʅ�`��Å5��� �"䌾}�����#<��G�� Cuʳ	)�$ul="%��c-�>,��q�۫~����!�I�2��O�!��Z'�*������%�66�H1!�$����Nx�u��}���k�'䋎���e/ �x�k�}� �@=����Ϛ��m���ƣ�k�����w>x��L��|��!�VD�V�#."�OcŖ	t��	�j�(m�|l��������$t��Ӝ9�'
�k��]bOt�>F/,��ҁf����'��2�zB����!0]��;��:{����y��ȌXq��ola�������9χ�4��x/�}!�����K��)����l��0�r�]|��P�*�]���+6�G���)(���a�2��	}��<�3��j�ל���|$E?̻���R����N��f-�{Vᷖ⸛��ɞ�:5Edx�E� !��D�%�lo/c��*}���Ed�S-�j�#
���UB�j\O~>��h���#�ʤ]U��[��@)�[`u��&Ӏ��������%��2�ŗ"R��נK����Τ�G�;ckr��⇎G�Gn �<��R���P�������ݠ�B�f�7C�����cƑh�(🜐���0�x�,ܰJ(�Dj�����5{�.�
@�(�Jl�0hHlX�,G4��蕵�����2��>��|4���)_�-.��+v:Z��-ǲ����(�/�
�d*�Eǎ������Is�^����ʬ�h�k�G���!�R���i�V"������Zdf�:�j)���:��y�q-Lw�DR�]�щk�?s3Wʁ���lMN�\����%�Ʈ>+&7���g.87k�-֖Xn���B���|m�/>��ӻ��� \�J���������ŕUuX�=��-�����)o�47���-o�1.g9P�x��3�9�b�}��V<;S�i~�.�LH���~%�շO��K�a뮯�L���̅���A�G��"�+1�+����KQ����V��nv>�^^@����n2M]��6�@���he����d�"�G�_�T�]9J�߆7�����ʺ�om���|j��F;�=Ԍ�JR��|���g���
5hk�+h�$g�IOI��z�\m��BF���t�|��P��]�K`�4D@�i
h����ŷ��$���G 2��J����TC �Π�ů�6t�>�^3���*K�#������_�্/�_�l���r�K����@Y�,��3��#D�l�L��g�Ǧ!�.�r�a��Ϡh���J�����8���L��k�T��3P��sZ�I�%D�BTJ����.�_������5c)�8{�{��a[��9���Aƅ�^h��XGd�܏B��o�J���xg@	ՠ7wEl8}+!<����s�oױ�'�}0l�N�ޔv���s�}'������ׯ�G�ry
 ��@���c���x˱�;��_US��LhE�f{u����;�q��w��}�7��������<�d�ڏ��7�Y
�)�N+��7�B)i�6��-�J^�7c�?���Y��Ƣq��
tK
��[� )Ն�)(S�8Oq��?kkB�9��2dh� ��*d1�Gԕn�^��g�)d�	hL@�5y��%�J��}���l&ps�� {��D=�IGN91y�T_�s�n-�q��R��SNF���(�](+�:PB���n��[J'a3�|1y)ׁ]U�M���,���fN���a##�<����7�ȕ���\?I9�|_U�/�9io �9������]ƥ���q�� Z���ӭa>%]���'���W��DGw
�� 2�����;���ʛ8w�ٿeJN-&��9C��-$t�,G\�sy�¯\K�^��F���<+3�t_��҅Z�_紈%�7	n怖GHg6���|��}����T����7Փ�r,��� mx����m�D	Rk�i���w>��2 �����t�sv����_��@���J]��
r����.�}]������~�[��I�<_8�H����'�M����~'��a���c�L�����=�"H=^��������f��Ùr���p4�(ed:t��d�u�Zߪ���]8�Ԯ�G7��1������;���@�/0 ������XQE�fm+ÅZ�E�#?�\��k�������&��̔��9O}�Qt���%,�+��2'6�ش��ާ��Z�_�����K����?>AK�)�qL��vQ
��</Z"��G:�j"q�UhBB�C%వgmc� :����L�1./jh0�p�o����R/i��!C&�(���*�]Qk�~��9A���九,e=�z	�����c�oP���`g_*��j����. (*d��3�V�I���SE?%����!��9�\��x�p1_-�3����Ocf�}��J���@��>��
���zg J����� ��C`4��t#�gг�e@����l9 F% ]' ��!1�+ݑn�3�e�^�����x?�a��9E~�(d˩�RH�G3>hb��?�]Z��m1��3��薻�f$�A�dW�2�0	-�]�ۉ���rA���"��5��P�t�������Xd�F5 �b;*�(6�@��{l�����	E� >4�˰5���n����V�f���"Nd�����1�[J��E����z�R�X���ۏ�p�/�,�Y�K�Q��3�z@�z�)zL��?�U��}a������2}��u5���˚�#���[n9N���7,r�y��� G�?���U��CS�߷ �M��.��&Z�D��[k<o��п1	�.�W�~m\^~�r��܎9ԧ�T?�x@B�HB����\��@#A��Yz<A����?���s���ޤ�ѵ��{�a�)�띒��=��y�OfKo=����[�S��A�*�6��;x���j@�.cc���rd�1�s��'���ݬLFF��8�vn;�A�������	�x'������.x�w����|�%�K]a��4�D��.�oJ�)��K���ne��������չp�\�R�Y�/
��^ ���|�?��,�l���1T�VP��,�	,�q��M)�d3Ǫ'���S�P��;���V
{@#���wCV-�_����kOC[[��B�p�PՓg���w�Ԏ��X2��r<�������t�����,6Y��oCm���I����f�^E���o�=�
�UxW����A���eOKr���$Ȝ�ﳴp��S�T�?V���9ZC\���;α渐m?SP�"{��?f�]�;�.%�9��Od`q�zH@���Z�2���H�hk�����5� S�"^K���hiG��C�6�
+��I�Ѵ�_��1�(�yCY'���3�a,��(G�ɘR����+(�?����DI��}�jcO���U͖yF��-��������ݥ�����)��̗��և���Wg�r�JHL��󵘹�g��J����Wu�I���?�������qt���T+���\������zr��%�y~���z�]v��x��煋�!CbL���r�;B�����x��<-��`Д���L5��s�������4��w�6O6rRvR�(�\�M��[K\񺤦�Y�Jq��s�Vz S#�r����I�*JIu�`��E�6s�X�"Q�f��֯]t�����o8ui�r�:��oI}%��%�������Ck����o~�OW��7���21��5�0��<<ĭ���ґF����x�w���7��V��9�|w�~z!�������u� }a��h�A_��vG]��+�B�/j�Wc����7M�&#%Q�w���f�m����1'W�s׾�jz%E5M��Mq�/]J�>/ȵ��@=O��0�UU�ڥ;܉�oI���M���t��V��gYOTy�w����nńgؿ���U���=dh���_HjU�C\^��z�P����'����lĪKr�!���CCk����k���@)�PD�\t#���݈tI#���f�����A��\�{?~���w�������<���,Ŭ�� ��E6j#��%E���m7�8"O��;گ+�Q:��Ȫ2�6Df�R�����^gS�O�U6�����f3�m)zfr)�=�;JT�sƉ�>���N�F��h�o�t�B���	���1�s���Q����|T�(A:�K��Y�F�r���1�8���Q��`���[���<�#�҄��G*/C}���qS6*h���`���2nP�Z��O�V�c"��NOSF��
H�?�:[�Npt����4M�5�+Xu
(H.�Qr|�Y��ĉ��V�`���bPg�������?�y��ؤ�Vs��B\���%nw��6�(x�[���B�TF��`�?g�
^Έ�,���3%3("���J���Kuf���,o�#���Ģ��r4��oq�%}[�#�+�����|�M�F�4�Թ|T�a����/8�&��7`-���x}J.�}�h�����؃���f��)q�{�}���*ܐzPǜ��3�R�p�C�)��-Ng�?��~Mu69�4�oFfP������[�A�}�&�?�6$����s��|�n���\�W��������sx���A9FI���6(���R�?{_��/��\�ӂD�nA?_ؤ��/�����fGZ|ޔ�uf��ݏ�f����"�El�۳�t�k���@q��'e��E�s�B����$&,���g}�xٌlI{�����JM����C���u�1I���|�:J5�ɧf>>���ļ�����}y��DGǳ��\Eai*"�����֕!d_�~�?k!�P�\_��?o��lz�	-w7�ٜ�-��t�;tj��� j�<���Hu��b�����jW�����@+H<މt3_�Fw��'I��?Cq�M۵A�||X6�-V���C$��2���{��VJq�N�<_6pq��
n??��Ζy���ks�>�.5�S��L<=5
|���ж�[1�bcU��"�����^��3������W�T���]�w[C7Jmo,q��	��-GQ�f�)n�]�J��OW���W�K��ҡ��Wa������U�^A�6�h�ѹ�	8������i��.Eףd9���i?���țN�i�l��'SJĝ::)���i�,�N8�TXp���,�����=��_��N�'���1�3�(�A��;�16���D�c���_O|�K��t���b��6#��\]�i�T�&���9t��Z'[���p�o�UO.����[���J})؋���3�bv�q�!~��-�x��G�	��c�h7Z��Z���`|�=c�D��F1Xeǹ�>��&�&�ưh�6�x1�\Z��gvj7�k�]�$�H'\���\:�M���������Eޤx��*гDe��f�g�����f����g��7�u�6�J����
	�Ƭ�I�R�"�d����w"��]-U��g���e�֊�C�"I�Tg��m���zn��r�H��qsfQ�au;Sh~�:�=��HF:�<�	}���E����\h�Q���%��ų[��z6x�_G�qjv/�;-�	
8O����∬�".��y~;Q�m3��t�a8u�.m��Ԯ�gD\ `��A�Vmvw�~�,�r`<�ct	L�9�8B�o6����p��}�5F?��$����㽵�6I�DF�(/�����wW����3�̈K�?���D5�G���f��2剢+&?�yu�d���փ^�ꅑ�G�E'w���/E��LB:��~k�q��(�L]�M��t]�g�j�S̈́�1�4w��[}Pl�L�T�J*��l��Rӊu�@B3ЪQ��^�t��u,��O5�M$n�2x����'��1J��R$��ur��r�U�M-SO����M��&ے�O���l��@���"2"���Np���ǐ��
޾�ǵ�0����wv�#�V%������=v�9�Y�y�j���*�p�?T΂շ��/���*	��R����"���?�C-}F��)A��Jo���L�b>{�wCd?E���j��f��K��pY�8�C�"��px�wT <)b���OuU�s��Q����e�TՔ�J�%m����)�P�h���Е$0>�?\��|m�&���s)�BE����86�Sf���j��А�1���c�$ؿ��F���e?1 >P�=Ղ�[f��>&z߷l����|��q뿐�Ro��ȷ"t����G��ݔ��ϷX����>����.����.����.����aߠ���w�?�@Ng! ������	��������ƪ����0K�Jcc�[��p�s���-�2�@ �L!�r��+11���a�/5W��,����Ё�
��ƗHV�ժ�vt��
**Lvm꒒�����6�9
��ʬ��Ȼ\ll{�M�%d�����k�Z��K���Yt�E����zVm���;?G�T5���\�Z{���h~y9�����]�lR����G��", @BK+��8��s$G(�t��Ѩ��P�DY~>d1�:AK��U�K.��U�U}$�
ӂ�g��<��<v|nn����i5���p�@�9�Z���+�-�cUFa�����h�G�͒*,���P-�ِDR�c��6׋��t}�:�P��W)��\�"m��c�u����3�e�E����^��Ơ$ats�\K���R�V[50FPz��6�����'��'�y%�$H����||d3���o����l;�#=%���G������\/�����|ae~[��f���%fl��N�qu�Z��@ꡡ>{�"��o��b�z�"t(M�m�~��e<�ネ���IK���|ڛ�s�oL����V�������tW�z�+�o�;�gԢz�Rv	W^�Au�t}CN��`��֡!N�]$��Q�R>����U-r~�`22����!&��kc~n#ô��-��C;��*�7f���ӭ(&~�o���)1��Ɠ��,�w���./�Q�7�	�����밌q�#�����Qf�a�˅�V��v�#������_L����^GD�Q���Cϖ��f{�b�+$��1<�����Ĳ5$��"�z``��(t;�>��
)���MF8�Џ�n�O�%�\Lk��	ߌ��k���TV#!�"q��Z���-�ðlE�<BX�Sc�jվZ}�M|��z��XnC�-��Y�՚�ݫ��Ý��a��PQ֙~�	�o�!͌*iN{
�!!��q��ߣ���-�u�X���%��
���'�		����Uvo����!��ټ{'Eʃ�N+۶�k�s|I�)��'��\#����k��}K���Dڼ����ڃI$,%�s>��qI�������@xnm|���\hO��1�?���,@4I�%44QT��Vq��%�Ҝ�l��q�
5�!�4�,`�IxO��y��jf�c��5&����'y���l>x����#�S�<!�3��LR�����褽x�H]�
���Nۗ�DH���G�9�
���Zh����uv�~,�A-�he�bHoc/\,õdڇɭ8��y�	M�Ί͏E+�.9 �0�$��$�c<'���-0~ga\�	���<��k$$�m�؛�8"��=]KEY�����qh����<1>N���;��Vhh(�R|�1��8��շ����7G1M�E4G1Ȧ��l���\uj��G�5��z��z�� ����%6�'M~�煼��v�����q���ut(��~,�~�&K��j}}}���� 
�t7������^hJ���F
�YWV�Z��	�������lَe��6)��0~�HcSӠ����x������?��ʃ��S�����/ۜ���?�ۿ�Z�[)�hɔ�^�?YX�ґ81�\�"������+	��=X_��lh�O��_�ǱO9�����rՏ����7/$ۊ>?:��p��i��@w?����T����N,	���'*_Y!s��������<��Y��3�?aD#+))Y4���!�h}Y��i��'V�;}�矍��!L�8/�bG��A��Ǐfg��1Ȃ***�MLccc�-,����ero<+/+�ECC�[����F��)��r2�z/�����&�Ze�6��>�(&�Sv8%x�$i�4Q�4}�N,����O[������-X���'�� �_���,�[�㑱��|%D�1
FY��p���x���U�(��񱱥e���h
a�4=l����H6ICMS�n���̹.�vHݕ"sK1d���G�S��-چ������;�q�P(�fp<���y��ő?������z�$))	}p������O�~ϲ�	`*6�;^	��V-��<��C��T���@�E��6
��c$2U���%���+{�;:O����Δ���x���=>nC	���q�����������3�����S&��^(������JE��)9��=�+:��y� gE��/�Qu��j������"G��*vyg�|���hp��:k������B���������=�LyO�1�����j���%�h@[���3b���n������$����*+E߽k�Ȯ�2Ih��`bbj��t���CĘ^қ�����RP���5r<1A&��� U��Z��������߿����Ϸ�sIn���2��Z�i��yxxL�aP���@�sc8=_�S33B�ǡ�>���)I399顷	�J�+��}�VQ/��Xd�7�@�"�#��Ǥ��5�Q ��s{���bw���i��술弹����n8�HԷoߪ<��+Pwf���WFT�+��o^ y�Y�x:�~�^�v�:>���
���������pp��LYM���-������r���g��{��E�^��JF�qWS���� Lv��ήA�������A fOK���!�kE�.��t���D��*�;.f�)����|�(��h���'�㍝��t����/�η~�^�ALBB��~�^�L0%�`}����+�8�-�����m����,)�dS�s�#���_��Z�98n�8�0�H���O�'��.kXvL����{����f����nVۚu�z9���'���;+wm��G��A�A?���H��v����n[��5bg�2�o�G�!Y}x&����r�j�����.S���8-;����+�k~&h�^XWOOO,�A�ĳ��������%���^Wf�<�Y�?9�������=o�O+-ewqqI������v`���_Td�R�����MѷQ��G~֌���8[��.:�Z��oً��3
o��#A2vWx%/8%�N|@�UY/�LWYSj��Шit5e ?��\Xr��[wF����A��c�3w{��`�X륟�2���5���|@�hz� }s����.p�����lSѿhʓ�IF�a��ؙ�L��zzz�c`����w`��,��okk�HIK�{�7��1�x��]^�<YI�����V
�H�*��{����������R���6HJG�٘��)C�NcCf��uz�l���7����8���3��M�y-���Y�Hn^#22rZc�@B��R������%)�v�f#'�L��o*:��:+U9�!Qe�쭬
P�P8=dX�܎�DAAIol�i�Y���6�����g��J��	�:#mO�?��ZR��.d�qJ�������+͍�Q__����Ӈ� =��'O4���Pvh_[��[�<i�N��Ǹ<�٬��7��RY����`�pQ��*Kǥ������Đ���\[��_����6�a#�Tu�!���OZ$paD�d�p��3���CҪG�)Y�,sin�dhd��`��5ⴟ���ψ�
�I�Yr��Z��Pv�?P?�0Ր���{j�7&+���nn����]3P���}u��t�w��zO:�n|�Λ�a+�iMNM��2�7555�l��Q��(�IK3H���&�c�_&��W�XKқ'�n��6���4����4c�X�� 8�^��J�������{z�ޒ�.��,ܮ�H�&:�Mȁ@�\s�H�0�78�B��xp?���P��/q Fd9R��[�չ�(cb��@�YE؍ɇ[�9?��h��S���W�YoCA���!���NT�{��N�S��;��,���.Z[�[��K��ᥘ��p= �ON:~��T�%�r1J���. e����2���˙��$]zH��+.���t;���c##�߿?�?~,,*�ANS�Y Bm��>i	�y��\ `'v�qi<$�/4���Ru׾)�����G���}������S���q�G���;yڻ��4ȆΥ^~Y����s:�`6�%�~Yu����B"�@�����хiG�Ң:�j�$�+C��A[���ggg_;l�کT��x�*�+j6�������x���IQO��>�k�gӌ�t�\w���8��$�5�Ud	T���<h}��Q���r92�V��>���:��ڿ#ȍ���|���F,��N���r�蘘��)�5�ܗP.��F==����_�-���og��#=�@���jrp�,w���ea�o��E6{��"�j��?��Òn�&_�r��W�l���B���@H��w���ӸQ.---τ����������̵r�����K�\I��_�l<$���z��7W|b(H�nkru{��@}���.� �H���p��n���v�N���z���KGkQ>�$��ܐ�)���%��\_53*� .� ��$}��'�� ��ϝ�ʷt�M>;�J�47����XѦ�t��c��ՃM9o��@M?����w`�f�˫B�z��ug �Aٍסk�z��H��`"m�g�2�h����~`Lv�;��u�@�4X����r I����;�'�nv穵�S��Ĵ��e�5� ����慔j3�Yt�R.����"���sZ��o��ܸE��7׀�$$&����_$ƫ�O@��4��1�`mOO�=���=�Eב�s��%���(A��;:�h�XJ%999 �b7�����s.$[ۉ2AY儎ix�����z��sr8}4�P����,�1.$�Ԥ�l�O%��"�:.�~w�H	��u>_w:��=c�����pM�Rk����E�NUi��ޚ4R���ζ<�O~`V(G������\(䗗]�H7���%Owy�9�l�9�N{�S]�F�xf���)�g���4�[%�%&ݑ�K�ŐJpV�Y
�J��ڳ�g�g�%|��m2��S��H�Y����o�5���2�\Cv���D-���؋j�2n';H�Ж�g�D�����3&�p���!G�^I�2�ׯ�|��L�IMEv�iN�yi]�o��.��HpEEŦ/ �Z6��3��� ���������>̶��A �=��C������V�40K�蘙������U��}��GGG7W[K.�	�otG��c�'�Ǝ�C��������݊�0����K���8��� q�a8��{�:!��3���9�zi�cq򣮎T$�Mb=ڱؼ������Lv���-�_k�p3� ��� Ʃb��yGY^锡�#:VVQ]]J�)���/��57~������wS�睋a��All��;IF��>a��ؓ�!�[4��Ett(���t��}��c��������'0 `�YU�ͬ�|��@/3�c%%�b��w3.��@���P?kp �mo��f��ؿ�XH3��B�p[a��H�r�Ӄ}R���H^B$e��P���8V�j��ao�+�'^y	Q��N�q� ���FH PMK�7�D�լ�u7~���?�܏�٩$���h��&C���?���W��Կ@����G&;X�:2b��y��w���S��eݼf:�ߡ���X�^Y]L��]f�P��Ibjj�56?Ӡ�({(pvV۩�bo����R��b�m�⷏(����"��EQYy���p��e ����S�'x�^{��['m����	���nV�o�p����v�P�mm����ѱ������^g�p�0�w֘�Yc�����zr����aFv�(=�'C>>>ՙ4��ǧ���:e�Vf@`�;�I��e-��rź-������P����ʆ���~�O�3lo|/����P���l,M�\%�*��\���jn^^DRܮ���I��ྏ��!�HU��Z�����,���x���z����R�f݁}rv&���Q՜�|Z�_��"������m*g!⏀�w�4��>`,���92ǘ�$�GUU���,fl\�{�ʴ��^����	866�@�3I��9w���C�TQ�_��^ZZ���}�g�&$!imjB����i�n_/�9�����UO���	Y[]e���G��}�z��
�����G�Sd{D��z�T�
]儧Ň��R+W�������b�]�!.>~ZII$J![���du������A-�V���M-���o�u'�?��������cv�668�lP򪄸X�YϠ��� �j�)�[ή.������N�DEDx��8�˓RP��||n��f4�O`��xubqQ^J�;��G��'�oٽ�Z��h=�7���&'}��W^N��Z�m�1?e���Vr���AV?..����b/�~�~ʢ�P�>2�1)���N�
66<�����륨]"t�q`?��x�F��tt䪃����/6S\=$*-�{�I~YS�Y�m5)~�c���B �ڞ�j�i����q�d�U�������C�U�*̴|�+��P:�hݎ[QI)����A�k��yyh,*K|���-d�g���@��#���]�A��R4Yjjj�+����!����v�a�n���wVx�7����M�����&�n`���ʚ��~���;�Ӫo!j�o��ިEZ��Ԭ�`y*DO#�\kk�`�B�܎��%+�j*��3��~O������I;]JD2�(R��WNɫ��GGG�=O��\��I��E��Fks�%�4X�0��L4{�ik謡adD$��\"�dj�

:yo�s�"��'�7< �N�3�;
��%�����C"*��֌���8�����$�(��?�y@�*��QQ>55�kv5 �)�؏�"���q9֏�\���'��M�]$P�,%de>�v���d"�Z�u������-�����wl����X�!Guq�i	%K�O\�4��;s[���2�r*u~�K~�1������]��'�;�%4��iƅ���OXL����.���y��Q��+̆��Q'�h7�Z������5��ԿM�&y�28�K�9 @L���q�`59��7J&��{���$��ށ�"�UW����\l�Y�����R���@�����{�N��U6�����de='mGd�Ӝ���� tMט<����\���^$�HF�W�EY~Q&,Iiix2��פ�ޅ����_�P�z�p_�p仳Ѹ�O�-0�	�� ߜ���z��LMǯ�{VWa�Sw��9������Io���[`�x���nJ���F����"e��2��ϰ <���V�X8�ÍVJK��ԃZ�=���|�p� ��ΤS�w:�v���ʛ��Y#��h��f�C��Rϗ����Q�L�+���]�O��=,�z �3,O>~t:8[����%��k�:�VU���/�*Ef��+�+�(*�[a�Is;c�E��؍�/������mN���?�҃=~ힹ�P�"����r���/GI	*�S�������(*�v
==}s_O��Fzlpڻ��!!�I1z��g�M���Q��ee�F$?y.!���)@�]�o�Ci:���&�/$���넅9�ͻ	�q[����!��j��t�����ձ������$��'�P��B����x&zkO�2T�d����Kr��0�
(��)
�Ʉ/%������iن~�w�շ㿼���3XX�F94��ڀ���� �0<�.�i��r�'?;;�u�@o����U��z����Tt\kTl��fAN��TTJLܤ��`�lB*�">��" t��"�#���ߧ���m2V«k��E��I&�Fvff�^��*>"����߭�E���w|/��t�9�?�"�"��ьATǅ|/�8L���K ��de�����?�:j0�C�o���P!:�7��Lp&?�^�7И�^���8���,�/�+���G�y��� O�:
��/�q� /^#�f332����A�����L_�����o�;�u(h|�t2�1��вa73`F�א=
�-�HK.�V�]�\�]Y�3�p����΁�^�4о ����K++z@�����F,�o���R��J��AH�hEޜ�����ݽ�\ġ�&&�3�6/���y�ƪZ3H�}!T���@�!U�c���{�D���x��ІGG�rs�Ƥ�S(��8�k������y��ꕘ��s�n/��yiq���	s�f�A��@ڋ�ⓒ�̟G\O�><J�b�H������<�%6jSIII�Q?9�h��Q~��-��Ю��OH�NO�g�gF.�g|�n��X,(�"����x�A��û�;L8�����wN�ML�͵ciBU��0:�2@�-��͠��)\�U�39�u��oԄy��w�bUmm庄A��*���E,8�}2'�I�ig��Z�B�rwD\������]]�e�[���(r<�q$S{2�DC��aVRE�x�@�w���ۀ1������%%��=o��O>fҭo�*�&(P&*�m�8!��^��&(x�����A��H���҇���ts����E�D�`�����歚�9Z�(�y��l��VSS���������(���ԝR)�8Ԓ�o������U>Y]]��R���\;"�������ǫ��u��f�4J6��(}����o�	��y#���ӺRC�b7N�]�4��@Z�02�m�K}��>�X�O��!_6J���A�t���766t��8B��gTp���~Kא7����}�,��ۀ�Zm	!n�//-}�� ��-�̅T ��6O�,�Bv�Z`;��x�V�E c�`��z�C�u��`�0�Z[2�k��B�#�7��.Z��"_���y8rX�nfn'����׷��r�|�������W�{�����<jt?VC���>Q��l��s7����������v�u�9�yed��06��8��-�99��z��Xw?~L�¢LI	@01�4�����
m�f"d 5���m�c;��W��C����o�#���)�4x�����rtt�e���$��Q�Ĉ�ls	��RL,rw��_���(b�|����7��==@�@�t?�|��=Lxw�?��M���g��Xcc�*.��6x ˜��Ѕ��� <X�FR??�R��o 4ʷ�VV d~VVƱ9SK��C��I�����dQ�oh(b}϶�����"�K^�o�m�;x
���5**]�eJ$%--
hU���f/u��H?jim�I�C�-' 	}8�R/��u���:/��J�A]�}U\n'��US�]7����@q��&y
�"53���1`QV�O����z������+w�w���%T��=��Tì��� �2=1h!��v T(�i9(�_�$G]]`��������/� x��zi�Bh����mT'�9�U>�$+S�7P
��`��o�C��9���?MT=���`��kޮ�R[�Fd=���:tKa'6ټ��d�b���T�O��up�����e����)@�Qk�ka�<@D��/M)g��P�D���s:�t����E��t�� T��
�J��pk:����ײn��E�\^Fx�G�d�y�ί��7@���J��#{�Ally�����3u��}������}�B~���@��sM�w�����z���@��xv�t ��Zd�5w��zba`h��5d!�u�-�xz㉴̏�>ߍ����g�X�����*������Q�z����T3B�z�z��(�Z3X%�BBTTA���/j4�V�D \�C ^IX��<�=���??a�|o����"�
����%�|�RymM1�p������z�s�TՈ��39��?m�4�Z{����@{�fjߥ��b�(q��d��%��"��_�8�8|�r��J)3(�����o����0:yα��s��K��D)��JWM-��OP�=3K�����=C�"..5��tɟ��J�?��W��ځ|��L������`�:/+S�������_GzLD�dk��>�9����;��������~��QC8�����H�<����f����a2b��6���(���D؈)�TY��L�D\��H�F�2��I��P�%�����!+�L��R �Q�U�z�*�E��ݺ�����|�~~�b����J :�>����"�7o$W�.�6�J���<][ۉ	/&jG;E_p�p�x����� ��z{{y��d����%*��U�-O_����`é����ٚ��@�Q�&ѹ��i�8�..� �4YTƧm,K�H��(!��Yp�b6�:��tZ���e���(�n�!ˏ��4�e��_gn� �����u��yfʭr=B�y�������y��Ey&\[|ܦ�
��Nq�H��쑠1����t&�>��ϟ?�=á�_RZ
��Cj��Y��`f�z���v�v/$ M0o�eފ�SUG$/Onr���F�Q`E��6~����V�USSCG�1��>��ty�6>�����3555�<1���)��F�Ё����-J��? [�����)uKC�����X���"M��tQ*�_W��+�Þ@������WUS����1��� ����K�[ºt�30�~�{�D5#�A�����l�X�y�o��	cc���Z�ݡV���6�b򈁛�{5؞n��/^�H	ޙu9V��˹j������T+�����	sU����#�!a��jC]��}���EC�:MA-1� �\O�}�u�G���dde�>7��C�pq�@��ֲ֝�Y��U�.��
ׇp�{xǿ�Xp���Z6e5��Ym±��D�uxu������#���hC%aGº�����8S�TB�[Wr�=:���Ti�D�����;�qT�����
���¾.�US!P�� ʋ{2���zӗ��a=!!!����m:����^���z0g�\�x��na>hN����K���/��_�
��W������W�j�@���J����Y�Tt���Y$��;�hh�JJ�BȀ���eggzs��A��TtL���3\�Jf!Ê�m����Z]���i�(���9��;����t�9��>�('��u����꼞�/ �$f���=��z��=Rb%!��`N>a�����@`^���K/Q���"�rƐ�G���sI	9�@���J%���xv�!4��b�T�2㥇@,nag2���r���6�Y�?+�����>�,�aKx��L�;���I��/ �j\w�0�f���S�/e����Ӛ��~�����5l�5Pk0�`~�g���{r����?@�SNN�_�X��@�:��7���o�UϷb��*�|��>L�lN#DM��RƂ�fd�_	9y����=�|��ja`d�WU�j"�	fI-򅶼�~ƚ�G�����̳����?B١���g�I7@�l����zq�p-�z
�����`��p�=����:��V�	q���"��#^�9��m��E�M�ň�]ja�
��>�J��<��۷��wl-n(�y�&me��0*��Ǎ �?�8�>V�v؞Ωr���@ԙ�5( `�,9�se����.�:ff%J�gy�/���um��I=���y3�!`I.�=z�������� шCE@��AA����yRؤ'��׋�@�������YY��E�c���X{����7��l�����pm�u"�o��#��RC�6:l��UѺ�Ǐ�����2��@����	Yo�����r�Dv]�{����;����x����j�A���v��@�f��{�xS��А\�� �E(1N�H���.	:C�n���Fp��y�5�}��>p+�	w���8���~Y�������'� T�@����fc,�x��}�n�s�����>��NA���^VWz��k�TXZ:55�����P��Nryp��}�j�@���Z҄�yh$sk~��%�	�� ���B�z;�bg��	����qrUS����&_qi�{F}����;j` ��<|�Y�kxun.��~����`_&�9W9$�3�?����y*=Q�@��m�3C�!{�%��I2�I<���*
Z����+�22s���� �*2O�������WtC�(N�ܬ�#UZ�}�^@�=�)\f��r��OX���wT�8������{�S[t��ti��6����5k�Q�KH�@ ��D���|&\�Pˊ��
h�(�	���7WA����u�#�>�����f�l7I	z�� T%6 ���m*���hd��r����,"2����rӄ�<%66���\_aA>:ɘi9vc7����:1�u��&Њ���G?A9��6�N^~�J�(|�=�n��˗r������w;R��z���> ��C|kC]]}�4h$�=��1o��T�Rޗ�=���J��`������:U�''�QL �=�����b�<l��|�?�<;^�ffTi_��_-.�`��� �ٖ�D���3`-�It���Rbj�犡�T.q
��r��QSzVV���$��ً��'"X��d�t�b�_@م���ql�ݷO#lFx� ��\y 
?

B=��1#�M�����p�e�1�+�Ҋ�х�����x�_o�k��Vp2���x�yi�Og�)i��@]�vR�2L{�A��+-p>�	n��;���Z
����O�=�`�L��KJJ
�N�O
����9cZ�<���s��	d�ǿg} ��)C�)JČ�+��mu�*��2MUyt���0�?g�ſ����E�	���^�<���(�{~>:�i���iM�͙<�i�j���x����ۢ�Rk$8�O�WB1��OE�ZPE�t��{�k!��ԏ�|EJ�Q��Qz��{h$�����$�>������;��耴�����iI�����"@O�Ԕ����'ȗ���f\�Kh�,)�	�!ʊ_BIBE�k��} �'�u)��	s�r [�ro���ޚ�*��	�=umm�����w��fZ[��� ����㵊�Fw�(�x�'Zv����x����$�/�GFF�N�KL�s���{ ��-�WN�t:q�p��
��ɯ��ZÍ����æ����PC�5���||dp8\w�N-E��/��.Okڑk��DwX�7o�0�Pհ���EgǻelҌ���~�X����"!1�������|��w���P��o�����$�fP遝�[/�	�~�^��a�L�h8�d���	6�<���W漴�(��[.&OGN�[ ��ME`뚲Z���x���<x���nQAAA.��c֌��_0�VI�'u8ܜ%�,ېO��H����0(�����_�^s ���sI��z��x&�f:��Ƞ� 0�𲆬���k4��S��
��NWO.���~;����>Ej�����(N$��\2{H0}��Ë��^��~c�wCU��;;;#��h4�����{����h輸4���j�AL^3�����p33�݋+�0U�^x�E���}�7"�7���+�M��\~æ)�.��s��[_�Nw��w��	�bG�Ƶ<|���/�����)��?�Ϲ�-���:mV�T���M#:%L:3:��c��E����n��A��lo���Ę��22�i+�}N���Dt��~�?�©f~a��D��������E���wO��wXӏc�y�t=�����3:&F���k,�c8}���@Z&7:�<^2����hB5ϭ$�s��u/�W�<_��ښ=b<(�����ᑑ���(][
�S$Td�>9���*H���N6^�C�ӏ��������	�//D\$�����-#�@;'4��{JNM-p}���]o�v�Y{���$���{��u�3��.��N��o��-�p[q4YbccK9���ꇈ,2��ސb� ��2�
X�;Ӂ��J�S����R�������)����c�a��^##JU3�-��dZ���QS�1�����&Ɵ\������	�^py���* ��	+�V��)��/d��A_W������K*��nZ���r�-�|��4Wۮ&aݥ���|~�4.��{/dm�gI�v���־�?*凗߾�a		AZ�Ŝs.m8�۴��������c!�S�k�&������De����Lp��p��?���~�P�ٙ33���N��N��>77*e��	�e�8�LGg��V1H���;����sk���_�^t4.�y_鮫g,zzz7����\ZLY4��� uww���#y�� �a�S猱Ќ�B�4�%W�"u�j}�#�¼k�b�.����i�����}�`Q�mt=<���<�F�$WT8	�(����HQ?{�{S��Ӱq�!H7)�"�x�����ǭ4/��-4d+�$P��4��#�j�oII�>n�ȿ���jMk���c�a)��:��ȃ_$7Onz(O�%�;5^�s;7~���l6.._��W��F?K܎��A�"y5��5���OS�����뤾�j��m��j�_����2�dM�EG0��5{9&�#7o��p'aHKK�2�`x,�]D��ɓ�?Z~����Ƿ��ZV&B����;0�Q~AA�1�͓n�lCCC�:�+���w�E��#>Isr��70������mn��KF�Ή�>	���Q��ځG{p��u�%�H��;�%��E��ԓ�`JJJ��\<F��%��Ή-?M���
dBK;ȳ��|* Ⓔ���TJ;;;�Gtu�JfdR�����%$"j��d �ch;��������y��(�v��㏀�cy�3�]�������T<P��UU��j��=��-�/""R�Pf�	�W�i�] ������+7��\d���M���0l����kb�Q4l�zB"��ji���������/^�+��)�GL)�mƻ��0�"U��#���f⫘�M_Z^E��-�0g�	�.--u���!��LF !v �B|�jz� ����gp$��֗��*s��O��4,�6< Ff��CB�)�*:�ZQI)'�����%-;%))	�����H9:��ڋ�U{0
d��uڍռqQ��CFO�����?��=6@�U��oE\p~֞?7�)IA|p/,q���_ �s����$$#���?4\PU�۾*JK7HI#�J�t#R���������K���p��n.�����ctu�=�>�{��6���(?!�Ȫ�X�Z�v�T?�v׵}����Ā|�D�\h�ˠй?�<e����@*��h���"G�����5��g�^e��1�h\Jj*��D 3a���
�	/ٟb �=���l��F����CY�=��
1d�@�Q�I�*=.nn��4>�aI�T�Oe���d��ie7[���{��1��j6++Tx����~?�F����kKy�o�'���<�dڃ�o�D�/����-1�.e�?��ȀI075��V����ݵ�^T�`u�[l�G�5՛�=�j����!5x;�=��u �K2�V?e���v����5P��*�LrRܸO��ǥyns�wq�FQQQMO/� b�?H*$$$V�IQ�b����+�#_�Ȳ�pe��g��0��ŏ����i;Wd��^���5�����p�kVo�"d��-I���������FG5��Z?���0����f�4ZorXwx$�a��C���4b�E�n��
�H4O�TQf��ly[�����
����8V�ԇ��Gȗ%`:���E�7e[PZo�26����Le�w����rk0��9�G��75E--�))+�x�↬4T�W�,�X��'~�:�a�J����#x�'���RWW��7o�n�Gl�tt�����z�Q	�7=���j����V
P�����п=� P[��gdt���:^��m�տ�gP�P������$�9���K�Y�x��]ͦ�A��`���3�G�������Ԑ��Mi[�"*�I���y�~���}���XN��꺒3�G~��<R5�[�Q3�}z6\�g�`��f����K6�w�+����n��IY}�b��W����6��ũ����DEc���|�B�������3�cޟ��p�Y6]�������$:�O�>@�66�+++賓����GU�����_N�ۥP2z�\I���%���h�X��[n�[nt<<π�W�ބI�/..�쟺������gAc06��p�+��}["�7�vr�%(yttD�j��<p,D�-\%�1���E�Y�Ik�r�A�Esomm-�~J)V�$Z(�5$��J_?�[L,ȩ ����^�L8���3��Ȉ]/���D^K�&r;�[��,A�̞��69��A!�R�<���I��-�;8\��&�T6�?w���dW��f&(AsVC����j�똸8s{{LoooR��3O�X93�qp"�`�#�1W8⡴�����L~ޗU.r�xxx��� �cB/�s������p�<�G��ݟU�`,�&ҷ���J��I�;��pv%K^�=��`��᫷oɶ����|�T�1Y��$i��v�~�s��"7�}�Ӈ͝��*�DZ�E˄IW9 �mmmM�Ξߏu.�v�+{�2d%��7wf��	�B;�:��^瑃ܮ��RVV6��j� 
����Ps����,��F�y����xVu(�G^�:��~���_�A�ɖ���:� N���G��j�#,8��!��v"L��^�~��ʚ;��(�3m����qT��l����ކq��܍��N`TQ����a���;
�U��b���������dѹ���ݥ�8]��y:�L�o@tQoU�@v���F����`h---z�g�X;;;^���*���+5�ה�H�.��7�r!�x�y3��e��C��a�����a��\݁߆��1�J?�����o�"E ���������5ɨ��:�x9��^��������.t��"�?U����;>9і�^�&�\`~��&(*�W�Ẍ́����ˡPP-�ˠ�����D�n�S�x�P��I  ���)�<l����~v>��{���=�ݩ��*�K$\MMM�)�}-��`:��w`V��n&��p�df���q>��|�H���R�������zY���J_ד{6WW�l=l(���� g���{bI$���_h�6t0>���)�^��n��01;.w�/�F�מ�`�.LYRZ�dE� x��
���ykK��8�#�v�ڴ��bw�N�#4�WP��j}ccY]]d��;A��>	�m|h����9���}"�81h�?[6��n��>Gn�OJz�U�������$������O�*82r3�0�9klK8����
�TKoY�#�0�;1�0/���2��&��TP:� �fnF�Y����[l����S��RD'�$����G��k<����u��gMa���!hI��

��DLP� 0���0�y���='���uCq#�zƧ��>;;s�PW$Q�N�i��i5�;�J��'tB�C��(�V|/�edeß|2��&����k�T�.6�m�/hC��gR@��5�Gn>��<���DnY��~O@D$���M���w3BB�J��Xx^W0��A�C��������^�d�T@�@T����3��f�N���N�I�!�J���q�%o|!��g~���d��f�d��U�����W������3��O�$nB*�@S��J��DYp�=IJ|ɛT��7�p�z�,��B�G����>(�m}���)lll�V�n�&��:���� |�@<������Ƶ��"\pxE	�|�D������ʣQC��XX$����mǨ�1���@�1[��������:L�����-~T`;�]+Mzik*���WKV�0���`�r~v1�ȶ�����d]c�x�:�i;���;-�#B�#T{�����m�����-^��7q&��XL�%�u_�#RLD�I�i������{�b����)���H��4�g�����T� ���.��=���}_���=9�ʢ؝�z�T1~~��"���������5L���xAH�ڜ��{д�<���?qdp�H�+�C��Hx4��F`S;�U����;�t�H��*;�휁��9ƛ7m� W�i�x�J��V��WԪ~02��5v��]�3I���[_�i�2(��������$p�M8���\v�K,y�$'��ǆ7���{�)
�qKdqq��%����}\�;�TZ�;~6��<Ƞ �m_�b�O)��#��l��ɟ?��&��[|k�A�� =��m�G�l�יm��8��{��vt"�xY�����p�#�`�����]Ҿ~���&m_������'-���5Q�����k�y��D�Ӻ$��ْ�/��+���h��X8-",(��ʭ�w%D�3Ӓ����ş*�'� �YXXd�3su����؊���y�E}�&!"2����҉Y�L�t���J����qsq5�p����J�ʬ�"��n#���Cx��e�����<����a�3�-4Cy�%&����ݘ�un���a�&���������E��P�ʺ���y_�2uiok��kx��M��5;��e���#�d��O�8�9�h.��ք�-�t��}ɛ��p�	' �UwO1�C����ʓ�`��47t]�<֕�����t����ɍ��D�1�K��(��A�ֶ���r���S�v��,?lS���έ�TXqw���+q�2��O���a.�hY�GVG���?~�hbd���S�c��(���.�X�gr���V_[{���f�����}Ȍ�r7�w�<��Cq�9��~�ךW�G�s���R,y��������ɥ����򨙾P���z	*�u�7�Қ��^���!��D�{�
z�z@Wc�Ax����H��S��أX,������8�R �,q��e�vO�\5w���^M�����_�� =�t��yyCy��ػw��**(�F�E�m�/cR������G�3�M1m��Eb�'k��A��R��º�����.\W��A����is]Q�%���`��ߤÇOt������VB�����ә��E�y��]�F�<=�tfa,���
������]�l~�C]���S���KA?䑫Ȁ��{�
7,2��$�x�?_ X��Ȍ$"&v��6��s-��~���eu-�d��{i'q�'���H5g�dR���U�Hhl�ML$����	��sh,1!!��@��[��b͢ʟ�U؆/(��=��v�d���/��~�ՠщ�b���[�j̡�o`��xo9R'�\.j�"?�72F �7�����E����=��l�f�ð�`�����IiCg���� |�;�QW���̏_<y�=�ۚ��WY�M':8܇poD睂����ʣ�S7�rB�bhQ�u�d��dd������¹[9M�)50j�0\>H �P�X�vU����f&*&�g8ȏ������ ���=���V񷢸�� ���G��!��spp��Po�Di�7E���� �����VWA�G�t�a�d��"��-���0�����_�Ze��W�-��'���S)G��G@���#�QB^g�xb���B"�
����ڻ����}�{�I�pr���Vu�y��+�tn�K�rQH<�X�?����/K��Jx�6a�+�+��@	tc�#_m��:9P���.ox��τߪ�}�$;;;?�۹F��a�pQI�;�6��7/v�z�d�b��=[s����z�����0�Z!�����)�G���%��Î�a�ɵ-]��Z�ih�Yk���
j98���2lcf� ���2!�Y�M�H0�VZ�E�奤��y���A���}��8����v��Cs�q�DU4�r�=�*���n�?_ER+���iL��?U��oۘ���f_�{QR���b�����w�r������[U�7�c�Q���sgd�l����΅~��%��~d�/(�}NG�RSS�QY[OȏwU[�����y[��}y�,���-n�� ��j�WQQ���,FGղ��-%922*���E���I�dIJ�aؾ6��\l��aH������|>�yE��g&�����A6�� g�(�`���i�u�u=�������!/����W���R�\����՟X5ʢ��Tj�,/�l���q�U s�'�C�yY������!*�D�#���mHH��6����^�[�=�p��N���@S�G�,�?�A��C�!�����6k�JVN�se��(
(��)��^���wE�2��B����>1�����0=���7W
��_��!��>>>�3���:��GO_�u򕃌`�||�p��l���1�c=9�۹]�������錿ԋ��'p�ih�*[�UUU���T��J*!�
>��x�e��kI*0�ԟ������Ioo��v���\��5%�����8�c�j
���K3�U�o(<z�H��0W/  �<~xkO�J��0�,,�����h��4��3Ԕ���zv\-�f]C���.bf����f�em-�����%����򖖖��h\{?���g1̸苃�<�s��u𝹹�i�����dip'B��UVc#Sr�@�h-�T��+h��� N�0~�L]t�h|8*�n������E�)h�rg���q�����W��������?���8 ��ݵ��)�:��x�k�Ve��C
`�M��3���G�=�c�o,�����Ur�)��@/N��ɗ{�W�������U�+!*ڢ�4Ր�`��|/��	n����[��/]�J�4����+:���xz�k�q2��J�1O�*_⭓��/F�}����-l�#�@feXQ�Z~م��r�������;�S��wO���CPAw�)�srr����6�gg�*����;�;��&���W���J���u�G�M�4���/���1���_�ѯ��3t6�nTV�W���<�k�����e�{�%��i)����-�j����_vDW�<�^h�����������K�'�7�7Q��>ZU�S�l5�� ��RuM�3Cz�>�`O4
}��xM���>0>E�����o���Ρ���X�̑?�Oǂ)���L�GZ03�P��1S5h���,-�\]G�p����:��͛li�jz�~��D�g��3��_�1T߳|����#�8��g'lbC�j�����յ�i���@���|��n;^XLjff�_���k0C����Fq��tu -)%o�����$6�E�(8/��g}��v�#�;
G�Uo����̋4�u����O���ݤ��)����*��	쟪��5�d�)�_�^Oo�S�	��كhȵ�ښr\����I�����s��**�La�_)))���X��<<�@���wl		gՋ�z�<F1g�yq���Oȶ���w�! �X׈���ǹ��z��+��?J|d;V���d���~�#�c�+�����m�K�C����%��{(��L֮	���j�g[���/��D_��>B����*�A*L�z{;ШM�K�G��YYy��r�Q��:je	�ijŌ��r����q����a�regF�����1E��z`jl��Tr�������p�7����Q�0V�����U�UY�9���פ^�Dz�N�ҲZ�F��W�l�i��fEH��P��v��^W}XSdN�0fE��^�M}G:b��y��_�'�1m8"����Ā)�ǄN�e*,�;�n����@UQlv�&���݂�W�P�n��0�o�%)��G�d��_DV̾[XP���v &&��2�9�v�z�u�)'�d0��m��v`���)5���V�԰X�p�[K��Rc_�E*~������ʡ��%���M�,�$��T�}Ђ�>>4�Q[?�:r!�t�]������w��6��xWS���sf���	'U���ł@��A��ׯ_�(tt.�=�|77��Œo�_m����)�j��t��K7G�~���\�l���K��V�	���ۍhD��֚(�5�\���Խ�c��c�����[^��<N�,���AiOc,�JNI�|��TaqwKR@Ψ!�� �=(�cʹ����T8N),,4FY@�!n>�j�"!��V|�M�f���P�6���Vd�@mʉ�{��Q�������[?%\<���׊T\�Dj�$ǜ���PaX�{>�\O4��VQNF����䤿�G�`�#�ϟ?����˒�֣&�dd�!h#��r6��ZZ(�}$l.y���:i�֍��o�vp��QQ�u�wI"\��5��>�l%q�r�w����n�L��Z���L�G��Þ��)p2��6�����A�w��^A$��oj
����50�<�
Y^6G���W���9Dd���rW�o�,h�������c�/.���{����I���g��1��Fk6�����
��:`�np�߬�i�DmǩwZ�s*�a�A.��틎�N��2j���Q*�~y[���X�8S��T�$ȑp��R�2/i��lDZ�W�&�Y��s�G��A6N�ҡ/�h���75��{ק����
��5�5TT`?%������}���a�W���"�MXDĤJ���l�f�n�	F������j�U��3Yi֩gZ3ۚ�-��[�	����_������Dɰ�c��"��,؞�� VuM<���ඳ�ϚkJ�}XEW�*,+�񱶶��{�۸���c��������&��ů�|�
�LLG&w��GM�g�6�;�y�p�D��QVF�c�|�ڇ}
"*��iU�0��i*��$ee���x�	]�1�ޞ������^���(U��I{9 �GDɵ{�g���vmo��?|ͭ�M�sꊷ3���N�^)�GE5N����S_����c 4)�k�������M5�$���+�b�IϤ-��gH|!9%e��AK�\���r#G�4�90��RF�6��:�#s-����-�m�>��V{fA�о���8��(U��}w��fI)���0�[x�s���E�/_ű:rX���᝝�.v�H��^r"��y~��ɰ���������[>Z�q������	U���|�|�����?�]��SP֗�����*�!�J/d:�׭Z<7R+�����Nӭ[����ik#�����;W^��{!P�j�����߿,��x���D��k����������ꩧ�-[-R<!~X���͹�A�N=�=����W��%#}]|�\3��zN��O����N����a-��g���/�ߠxxYoA��>��Ņl�mc٘��aE�<�D[;��S23����M�S�Z7��h���}�wI��@^|�(�>��z�E��KXx{�UI�
�è)��n"I�����ݏ'�Ţ��5D�Ҹ��3@̇�w[�-WFN<Ol,�����]<|a7?�I2U�&����&�ĩ322(.Ex��*VBp���*�u�g"�GY.�q��7���	�L9����:,,�WzW�є"z0�]�DbF��f�g�w�Z���~M���p�gD�JKq���Q@pp��QE��^;y��:�~*͝��vˏY0����҇��ez7Pb��T�g��'�m��7\�C�b�Ɨ�!8�!lo���u+m��Z�s^E����ߐT�Þ�`��|W_k.��>��\I�Gt��EG�g�)%ԏ���>���7��o�����'eT(�wm�����ZY�����A���_	0)��%�&;;R22���Q!L�ڄ��o�̓!Dm0eu�t������(8�D�`>���
2!	h(^U��[�+�3��FS�#��p=�}�[�o�ў�s�g!A��4�H� �s:�+`*:��2��$�7Ե��� ��@G���Җ11���U��B6t�����{|r��P��F��x�d�o��K�IH�Խ�#8?���2X~Xf>�2E�7h��<�]g%==+�����I���R����J%H���u-؋����&Jj�<港e�J�X�jq�6����61�b,�cn���|p7v���8�_+��t����v.i��.~!�a�<6�j��;㖳d���[(jl�����鏩��b��l�����B%ڥ��!吷�&;r�ލ+&���,~�<�X�!��6y����b3���n��ؤ�ސ�߰v53Z ��^�o�t��ْ��wgZ0�.��gv���3�[o��i
����{\j��#�F�w(c�C~��eT쐐��C%xZ�f�mAu>���j�Cnߨ�v��P
q�b�WW���>�k��W�R��������>/�#�7̙q��U���{ji�/^\ �~�����_���9�B�'�??xu��̼L�K-i�a���V���Ts��aģ�~��Wt �8����H��/� �NXI��*z�K�4���}o_7�bUw�㢢��h\�#j�~X=.�ZҢ�ݖ���ݰ���(v}�*3/�������/	"��E0'��6�c�X�����c'���5?���Sd	s���Yj>��e~�،b��A��4f�"����9.�ᐮ�vX�
r�WI�|��<c��='Q�ѐ6f�<���=��3���X�_䕃�N�ӡ�:lmVC'K�3N�L4�-�L&,,,��;:�/DB��=n���S��n���KHM������@FZ�ϛ]���J,<n6���Xr`榸�l�%ѥ���4�����X��c��7�r�Aq�#¥"F�E�Y�DLշ9�����F~`��z:hSU	u7
�QSsbRׯp��yG'@݊���vtT�ͨ�_���;���&�Uq�nOr&	����g+��R9Zs+������d�m�D�7U�$�*)+�����Ω}e "]p�]x{�{��6�����kk'�|^�TVJzbk�W��_����5�79Q�*3��(h��A�˫��9랗��m;Y/޵]�fҙ�>{Ȕ��l��z��e�ZZ��焁����V׎��DR��Ƌ�ˁ�nY99nq�O�06]˓7���Q�,H�M�*�E8�Z�@����77G�����[[kj�T���s���Ԑ�Z/�B�em������s��C1��Z��S#��n�e_�H/��%��1�t)ZFL:�O4���}��X�zŐ�<(�P���[*��%�\[���Q
��#��@HG��=�YJ2i�������5��+%%�5�TLM^G�����G�fW>�T�#��zxof�a��I������G�\�h
�h��&�ж},]Z�Υ�q?	��B�+ .�Cڨ���0&(7>�J�P��VI���� ���z���=��6������y���p&_=�C�@�pE~�J�M����Н������Z\�c�j[>nn����&GgkR�����}���2R'�2# "B��� �&6>��������l�4)[79�x��NEwx���7կ_/w��C̔�	���U���~W[EV��ϙ3���Tcn}w�%%�Yb������be��Q/�́؉�%Xj)�;���y�G�M�>0��||�������Ю����4\\\AoR9H?���?�������aq���9���ZI���*K��F��ҕ����כ	T�q��!�	!m����FFF?���n����褰*�J�5ũq��I�(z`��K������9Þ�9����s9܌����:::�pv1�ǔ��]h3p(ڣ�����T_K�<eB���/��e���R-�P=��9;+�7SO��]9�r�)<�J,
$��p~�Vc�F^^��3�3���?/Un/�E��?r�Ƭo��FPu��8�h�-�JA�����ndz:��IX:_=T����\R3:�Cf66iKK�����>	�P��T]� ��߀&F�GAڸ�E�Oa����a7́�k�
?��w��be �El��	��s��?m�JA��uXq�%A%�ma�I$~xCJW75��J�r��$7ҝ�D�N�4�N�I���X��qp���~�+v������aLF ƫ1^�Q���KsE�I1�I��j����$f.�Æ��q�TZZ*���"-��ȋ�����)-ljd�j8����d}�r�w9cۓ�(dx�u�q����D�{����,>`U�A�� � #�6�WZ��˗/ߪ����� � ��[��Th�khHFA��M/��MF8p���}�����P
�d�%�������-�\p���Wt	�n���_]����{s�#��;UQ�a�j쳵L�Ճٜ��qKJJ(<ѝ����[CM�߾]�?�
���
� k9/�����$$Į������׉����y#�����]`�e�)z4AoRM�5"]7�)	Y�K�7^;v-��}II�&H���	��Ļ�*v��k������%<�Ӎ���;� �1䊆��eA�+q|_H�5t��_ث��t��w�f��ݭ�~�}{��G8���ެ,
䩐����%AɎONr�6ra�负��B@Q������-9�H�+))���q�����K<�W�|f\D�ۣ:��D��x�_�A�9nw��^Y�=�&~w�&������m�j�[��a�(+"��9x�4����4٤�n[-ǵм��^��#/5`YRR�xyyi(������G�����J��� ���g��qQhkE*'��l+�>OeǨ��>}���n�)}ҵk�
~&�]\t���b�b���Ė�;ԏ���׮	X��O�9��+Ϡ�������&�ąVB��O��LL����A�<��p(?�X�s���Qy����7Dd�H�?�B'�wX& Ņ)#��c�VS=��ֶq��Gy^��抝�r 
S�����hM��vq�*�a��;�vBB¸O���ڱό9�ů	��L��sp|�H���	���2�50P76�3��w�����VV'O���@u8��PE�m�ػ�Ra�u�Ŋ�()-���JT���iEcc�?�� �@fǻۋ�6�W+�g^�����jj����W���i��6��Q,�M)��zm��V��r�b�AX{����Ʃ������ܔFLlR^3���_�0����/J2�לQU��a��wz&���G�w�����>�5�_�0�!��y�d�Đ����O����G(��~���YfC�0�s5���YY����Y[��ф���'iy<��U�л���_A~�n��H�>cJ\�C��1�Jv(O�g��,{ێ)�ˋ�?9N�wa�Zڷd8xi�ȀAh|�j��,!�"�Oumm7ww��m�l�Oj������<ϖ�9��o�w�yT6��b����U�È��f��p�yU�����y�G"gT�Rs�N=i3�-3sv�Y��
�3ss��k���nG�=�͞���#ќ0//@�䡸�YKa>���}���r�X,���_��݊�g��r!��_�41Y�A��Օ����_���y�Z�ݭ߽��9"Vl+82�1M"�X�!-8���}�_��׵����������\g9;8Hl�,xWu>�ts�oi�G����aI��KxuĆVX;���u�3;�Y���ڞ�g`�pT�-8Z�G�vD�.S$h���f�m @b�b���3��[����m���Uf� _X��f3Bg`��7Wj��~_	\|�z��~�̓@�;Ȯ�˨�����5����Å�i����Znp��*��\!6�'���H'��u0CW� �O�9(�ku����4�&&1�,{�N/��(͢o��b�UB�%�=�R��|�l���_�w�~_�����$�p0�z�e�E���Ϋ�Q� �#Qh62�%�4ՔVz"��8r鯮ȡ�z��O@<���z����>ɯ������"�"%��TTH����tSs�����w%+j�ql�y�Edb?������r��ZS�_⮟����Գ@�޴�[P,����-?qj�q��A��m��yc�b.���Ӿ_�Q<�a�Ů��V��))����.��>��lW�[^�Cr~��D�7@T,��}����`��WsI2��F5�#�C��$�ŋ�X6�*=7�|�Y0V*.��hw^^_�O�וj�0t%98��5�\��9��-O�:�NY{�����F�6θ1�866�a�nFMWW`%���Tg�$�D�[�f�5�4{��+C	�����R-�	?����z���%�{����`:I�='����I�L�T�����:ۜms[#`CCC=��*��� �>�2RQ���S^�WX��k� X�q
x��ظ�cf�/��k(3ƻUџ�(��Tzɢ�ݱ�e<�z� �z��O��-j+%�.�v���c�T�k�:|�<�(^Տܿ��0���"����p���^0�c��?8|X��Ҿ��͘�=Q8����^� n[�X��>(�,ָb��4�������<�����]W���&
�e��VV/q�YM梀�1i0�]K��/M8�,�D�869��7�E�(��z����G�T����k\���|���j��\{�wH!�w�� f3៿�����ŅB�cbHP)��q?��/�ѥ�ݔ�����xW���w���@ʓ.ȳ(j|�ۓY��'���ߎ��ntS�bR;�9��*Ɋuw��hIM��Yx��lnzu�g<^MR�z&y�pu��ߗ�'�L����򳼽(����[��UZ]��r�6*�v�G�c��K�e��a<�&��U��9���Oƒ�0�T�������s����n��h,��(� �a;M����(>��}�^#� ��Gσƙ�pQ`��׭��؜~��ڼ�	plu��YQ�;��࿪)S��Y�⒐�(%{���8ZY�9���>�ݙ*���M�H06?>����m;����h2�7stՅ��O������~��v����K��Ʀ�7�ܺ�,��bN����4��dD�\8����<fUǹ&�l[1���8a����,!� ��Gj9F��Ue��6ic��dr��s;N����l{X������%��2���	����&���vD�E<]z��0�u�ں�ұX޻�
��|�LW��Y��S�R!Q�t��a,��Ǉ3��5t|��}ǒX�"�p�{(#�EȊ$@9e�C�H�z±��^��Sz.~m>�#!�˨��Y�Й-���m6x��a"�Q�r�Bh��wb�����U�ߵ��B�Ѕ^὆�q@���U��{����Ӵ� 	�u�����4��§��Z��?=c���I�}�?�1��=..��������^�P�@|v�z�{|*���dΕ�D����߸��ɭq466�
��S���T�l��ip=��Cs�`c��Q��1 )�B�Ʃ*9�d����3-��M��9�T���My�CC�.�]�c��ia����}P�o�j�zqݷ�n5>��o�9������R�B�B�t����		����B��蜱�)�����lX�<��� ����H5f�V_�w:`�5r��G9%%���{-u�`��Ǆ<��­6x�wWp��5�k6_#^o+��KF������`��Vo����g ]C�q�����1�<�� ZORP�m&��j?�*��ݎ|�5D�Շ0���`���ŁN:'f�05��f����M*�������SXD��]A܈�����_!KĚdzIo��KA���R�~.j���фX�t$OF��\fG����@�-�u�I�p������||�W��@lc������t.���-��B�j���$�LL�^��-K��S욃%c�B�Q��
��U/��jI��]F����Gˁ�+� �;�R���Wı�+J�=	�EdqҸ�şU%��a�M����{7�sX2Rjk)�3�(ۮ�jSg�%,����~u-_��ЃA˗��}��}y�e���(�<����#�pY��e�s��M��N�mM��"���ܣ�d{�!���w�������H�'r���YD-��҇��;��NMSs���1یp��l��ݧ�Ka�,��N�4�R?��^ј�0���jP�����.Z�Ș�iլ��)��vþ��t�~?�|W��g �|��1-
9y���1�<�b�b9��v��O�f�MQ(_���m<�J�W�зriQj��O��Ed��rtA�8��v��z.�H�}�����C�K�������O�6/Xx0s0O^/�NLX��SB��a�K0*�������o��G��=��[�������b�?Y*p�s�r��mG������+�v���w�Ɲ+���$�f�ۑf����M ����>[|�A�B���RAÝ������v�V3�[��<nC�Nu)��m�rYi���c�:!�&乼`����W�+���C���y*p�A#-m>1ȶ����U��}0�+	�u3ː�d�����@ގ�sI�i�1������������+��^��f��}G����ZZ����P�K��wTBn`�MA�Gݝ�Z��]�����q
��ɓ��Hv����c���l�b_ڬ��:�����|n�嵯5bC�D�W�%�x�M����*p]I'u��g�**y�a/�����Z�����0��In�ž��t$ddմy�OQCV�5�P�Oֺ�t�ŋ�<w{�gl����5�,��&��@ )�
4�k�����{r���H cSE&_|k3pG�89+It#�{upYQQ_�gG����e�Le�h�i�c#��eF�D��K6L�ȣ?�Һ�~�[<��~-`"1l5b�~P�&�mkU�hg�g�S �2SSOq��$8n�2�v��x�⿬��`\�щ�$3A�t���3�	-
�a$��׹�������[9�<Z_�(����:X��[@�_�馕�}ɽԸ�5��Er�t>�ut�p��NNN>21�8纒��T}�F�)C��C��\�0��Q�%���Z�� H�W-L4ekeJ��2P&7�EH�4�#����a����>��ɬ��*�U�&�)�����8�
���{$mQQR�tozJ��9�"*�kI^U{�:�aB!�a�p/D�r+�=3���Ǖ����3�^����,�>���$`�M��b����+���T+__n>K��� �*a"�H���gAK��c�1�9X��雒�@8�Vuҗ��m�hjk���&d�ƈG����&ߊ���^��HF�ފo0kKR�W�޽��8����IM��WWD�EQt�?�������%��l�͍_�qkFK�<QOO�^�{��x�wKxn�#�/eIi'�y��ϱyN͌���B���	�j�ͥ�������*M�^-��N�|�rk�@�Әm���UK[��W����Ι���a������[� %��4�c��H�*�J�vU�5���hw7�,ȡ����ܜ|����U����罎(<�!ф�^{Ur	t�چ�o��)� �£�K�����mkD~���i���x�ﶷ�f��'��fM�������LJ^g��ࠢ�j[�\\�vjJ�9��w+��V�WU�D�Pӆo����������{��I3��f-��+�w&��L�IH���xYՕ1�?�|3�5��G�s!6��}Վ���0v��q��ꚭ�8����l�q��n�ZR���Ũ�<��I&܍�_vm��R�]5)T���*��ۜ���<h��s��{{\��G7��4�ex5���C��93j�m��/�����)��9��T&��ʐ�M��e����{)�As�]�Z!az�VRb>Um	��2�<��O+��2�G�������5�y`���u�%�U�$E�䜜��U�(j��$�ɐ4�K����K폂��`t��l�w�R�
\��x���i���J�#c��s�@W��!W�֓Ehy\��F�8(�6,�E2�Wrf�C��c���y#�)l��&/؋[ZD���>�Ge�^M[��b��r�E%(�R��Dc� ��]���b�K~x����S��� *�	�$Q�㱢R�s�p[{����R�ŋ�%$��.}zf���A��sGsN���Y�E��& ff�2�(���rߵ�f����y�n��?�߅��/��5�NqI��g�'��o� {{{���2�3�T*�^�y���%8���hZ��5�V�l�RQ�#�Gm`� k}�N����{h�j�׫y�\��5z�Q;泐'a��-�yT�TUፏ����ͼ=�:^#���
����*g�g)�S�oon
� ��l��`��M_�����
"Hwww�,��%��!����]��-�J#���{��}r]�Ù繟;�������]�wJp{��!~0�{a6`�0���m���q�H;s����x��6�_r�Md�ah�8FGE)����qTU�(.�wYm�����k\�ap۸]���9�{�+&�7f���5�h����i����,)�ۋ^k��R����i���NX$g����	�!��m�^��c�1��}dw~�zdOV��RHH�U�I��88�MM�)m�T} ��>ݼ��s~�>=�mњ���_׈���"��:�S���	�� �Ư�߳�����:�/�c���$���U�Yq���!�Җ)d����%4l7[e���u������@��ڑC&NwC�]LLLK����hn��7��B8cbv혙�k�{
������v��V�xQ�9	P�>�R;�?8`A�E�	�hv�'��(�5nw5j>��HK&�(2�[Ո�bLZ�l}m�MC�KR�(�� 3�b?���l o�Y�BS��K�7�����nN�U\�= �ӿ=��K�2�#?���:[,JkcuތP��f�tj�m���.�yz�!e;ꙃ�K}����j�zt������%�Z������N\\(�g0���.��h�8ت8(I�����C�6���0�3��b�y��J5�"�2{�
M4�("9rOScdd��s��n6�w���V
�)���%D�Y����kd�>`�Y����s�*U�2<�#��B��@�d$q��^�i��ʥ�����h��E�	�Vm�N>���@�%,,J�-�@���D�j���|�0{�>C�O"��gd�y�O�\	��;�������e4N9��21q�v��G����-{C��/m��������Q.��Y`u�x�Ӵ�(��o�h&���cc��|�3��Zg�ߋ��̤W����Fk3�
�|ii�𝽎��Q�[X 0F{��	-/���֩jڐ��6f�b�n76y0癫'����-YQ�����8�1�%���0���t�)0�ɾ�0R��חd�f��F��c�5�����]��/���C�fs~PI����?w�w�(Oۙ�ꡩ�}}�ł�� ������ɤb�H?'D�|��(�Sn��*3��q��Yc�#2*/|��Ѭ�tAj!��#�2��ɰ�_F��D��;�)�u�RQE_os*0�:jf�%��%]9��p��۷px<�3�����&C����ݡ�'����L���/���[���wx�G�]lN.��j&s`q"�|�l��h�5�-�^��,��t.f�K��֝�N��.f�`��<zzz���Pqqx>�������r���s��M�Ge�Mj�����v�� |yݧ�_i�6�ڐ����[��e6�L'*��b�~��9$N�ع�0Ѐ��Wf�
���U|�n���`�P�o�-
�R��x�Ƚl᷊V��z�G��g�
��G�Hn}/n�V���5N)�s���|D����׷&�{e���T��% :�������D�`����L���)HSJ��&��4-ߘ$Qo��>N�Ih�Po༶_k�~��ۃ�~2X${8,_������,�a{rv(��?bAu���a��.�~[��(V-�����RR��^�ݥ 9��QE�=�H�8m�CЏ�=�g�?�΄w�#455�(i��3Оɧ2���\o�;�e��K�)�ZS�h���(}����9f`�����0���b�e��v��L~ssj5}kF!�N�;�]��a$�Of�r�T�ukE�8j���TI�������>��N��y���
ו}��V�fW0���e��/O��9~���������(КU�Sk�Xg�H]f�d� �?�k����7�g`=�f$��Ņh�R<_o��m4=ž�c���>���do�\�3Q�+W§]�����Z�h1�SX@K�ꁛz��\�`�!={���>e�. -������5�����p��c��b&�s; �aaa{]Pă�Pg��o_�i�G�_\�z���Ej<� �a�.�<}p�A���ѵ��;�5ѭo��b��^V�'��!N�) �1�,��U�z/;��4��7
o����{��s�؝��ۯ�*�w/���E���c'M��w����m{�킞�&5���Kq��Y/�ئf��J�֜�c��N��m*o֘�[f��BRRZ'���A�z���G�j]�v�ج�B�o�ߒ�>��pqŷ|�geRi�{#]��|���tٖCB�rLŋ�'U�W(�x�5�~�x@��3`^�����@�Fܺ�s9��Ѐq'�3�\jcMEp���׆��S�`�t:S���P4��Q�?;B�3�@ǡ��� b�x�DRD�����]�����Bؤ����m����5�=�n*��3�g3QIUdU㑒�Pf�λ�n0����F�_R�Zme{�dz����Q��J����!MD(ۑ���D <��� H��&�=��_���zEȴL���嬍��5�����h᪠����$�:�#��Q�Ph�������C���{@�U+̓pD2�^����v̝���V����Su$�/냜�sT��8u�~�8�:�L�L�[,Qr�	5��8rL�ʁ�R~K4�fZ�;��Vٺ?�����w*���&k�ח��*��b��'�,�e��i;�bBaK�л�Ku=��I���S�lI�<l��k�TD�%2fO8�+�-y��Xە����G���,4.f��ei,C�v������H��v�5j
_�e��x��Ec��100x��z�	>w~��WDh�5	N�7�i���#��lrZ�����B�FVG�ߥ�lpqp'W~�E�0S�1�wZ�lcpA�'\|>=,��������h|��膻����뚃�j�)!8̿�6���Z��
*��'��7���L�>�߁=�?9��]F/�i��k_])���1�qk[[
�L�v�"������9>�<�݇^���i�������l��$�UID�րO&�;��b��B=�MMM����D��0v����e���c��h�'����:�3��5z�h]���U�:�V��&k�p�,����*+��<+qs/���#A㛰�C�w�uŏh�k>��H�x��?���r�quu����;�<�t�:P������%��7WC&q+s��VC*���3��k+�PUi�)��9���v�����"�ƃ�݆�i���2�f����~u$�m�\̺�;?��~K����µ�y؏�:p��H����QuO������j<|z��L��_���륍�6��R���r����D�!v=滠��ۯe�g�2F|�h��̾y��))&���RY""�^��HQ(ss�M�#vr�泇����FU�������p�<Y�AVG����g�a�Z���\�$��,�F�E�%�;�o�6:���o��SXU�����~��Q�?�p�����O��?B��D��7���-�*�x��M6{�����a�����a�������*����N�E^�;�>d��p2a�F}j[/c�&���<::*���>2�@����P1�+�ˢ4�q�d_밂�"��R�3��pV�E`.�&):�
����b�w�������8�`�H�/�����)���Qs.���G:�J��
;��4���B6��i����0	*Bv����r��۴�M��K����--�+l�-x�Y���
 b]�-���7���t0��=�n����>���PAa�3j�EN�h���?��tN����s����{�����u9yy�M8L75�Cob�x��BMw9���/�G��1p�K�b�2#�>>VS��ǭ	���r���SRz36�}h�7��v8�+��A����|�t�ds=�Ã䳾�H⟡���������l��Ќ.k�6TTD�[q��<j��,[9t�u$�CC�3q��Y����8��v�)��P�˰��OY�4ޱ�v��VVʍI��i���tǢ_3���Q�u�^2M7�Dyxx�_bnFM����ң>��}��vkz�|�
 ,�-͔�ZQmou��oUIS���E�?}_.C�t�7D$��˲��W�dw�ӭ� ���S [�mr)Nz�^	�gV;���U��}�sl����(�zA��� o�Po�P�k�A��������Xe��S岍����Y�0k�qdˎ�c���1� Z���5ǡ�k��u�x�#nE;��aC�~�(&|�K#-m*�#�_���r�����WvS9� �	eJ�M����E�)�MMb����s����H.�;s#����y$^q�@�9�
r7��ꍘp(7�t]q�v9wS�4��mث��Tw���%\eT�5��%��o>�?��.s�-rPC3�F[Vzѐ�˄7��kb�\Q����ؘ}�ԛ-g<�B���"�^\��Cso�|�4(b ^ݰ���jT����"4��Ν�&��g�+h�D�%�"pD�<�L��]S2ҹT�H����H�7�vy��*�H�㤊�]9oP�`�5ȍR�����Ҩ>f�.3�3���6� I�^Tқ-C�e:�<�(pz ��{Q�8g�ۈ�h���uPa�r=�9`YX�7����g�xW��:��R�eB���=����j+�z�HN��\~��>���L� 䰸��s����9��0���M�P��`B�r�ʶai0	Y��W)�#*#��D���Iʓ�<�W�9�5Ct�'��;k����;;����vhx�pm�@LV�C���<���
��blP~�}Ž����{l,��0���Չnm�V?�ƪ��R�zZ��!�T4�Va��j6��E����g���_ODNv{�t�S����zQ�g,�.�!A��U��e��5j�+F�Mޚ@����8��\���	1 �u��:��|�S��ad�wۏN&C�*^�4�b,��@�v�ȝi�ڌ"e�ͅ/���ȱ1��%���l�n��0k/;Ftd�5��%①�=��-��|�jȽ����j厃�z	��x�����
�e��\����Tfn��US�:A:J�(��:~��D 7�N��-���2ω��T�N��D8]O"	10Q�b��~{�EK��(W2�!���U�����_�%g����P�~_����w8o�FM��ޕk�������9�y�*K�n/�����<�6|���_��ϯ	�	��-� �~�p[
y�5�;%��Q�*CRx�g��?���	.}?�`�6��Oo���̺1b�J�x9�6N�	[��lTYn�5�-k�� F��_�+���@8�k_���p��n�Ø����KM!͡���K��⚦%�H���K�4|�.Y��,ML�;�jQ��2*�d�e[�L41�hj�`l�.1,'���4zl�ÿ�i�sP�!��6?o���p���5z����1n�4B��j��۫!@o
Mk<r��Y��6�陘��=�5/�mX��w\l�I��EeJ��픘J9��[�m�DP��O�-�����ts���핟i�(Ù$I8-v�l���{5T&�P
��"]v������9n�^�F)&���?+�G��?X]!�>��Vi���k�̢�B�edD>ή2$ ��$��-K��1�j����{#g�Kj���ʅ��LRS�7m�x~�c� �IՓ�6N&�sp�(B�(T��>��Rn?L���xG����65��7��bO��Bg�	�m~"n)b��|%�DDȸ�܁�,9՟G6��׶����	2`%���m-^�F�qn	�����'q�l��~�lE����!�.Y�2���pYn壩y�����x�䚈��	3I[ق�?(�)C�+��6�
Kc�U������oz���Դ~����x�4a�sŊ��E���0K>"�ҩE�:!�T�� ��T�{j>�z������M�{�_��	��ȠG0�AP22"�cs.h�s
�<1Td�Cl�#?6��+�1y�[ݓ�~��}���1�y��UOf]���W����>���W�G,k�C�Լ��.)<�s�B?X��<�e�H�4 ���FF����� O���X�0v���b�8�]�M�/UW�����o�j�7^}�K۪�\ZQ�{Kh�p����Uu��'�2�mzkL]G�Ӹ��m�D��d ��*�䏗^��S�����&`��Y�����i���<9,�>0����F)�]����mSI��k��m����m�L���dcg���@O�P(k@��� ���;W&��ݡO�9��ECz���Y���F��A^�k���z�U0J�?����6NvQ������M�b7�@L��+.�3����m�ђtҸ�㺦$<�SEtf�FpDU6�v�l*���e��-.����,�J�dPy,�h�Թ��k_N\�=&k�3�W9�χ���W�Bh�CWސ����3)����S�FoCKQ0�ǙgG��Ŧ���KJ��v�f�544�<�&�@�s{���NΦa��ww���1@tYc�	��yK�W�8]M��]� �tFlB]_x�A�[ʄ��m��px7�<��#��ɱ�X!n�Q%j���e���,b���dz�sA��ؗ1��|Rr��������O���1w��Pm�>n
�@�P�;"Ƣ��K�O�n%bۙ�?��\;s� �=��w�4���cat~�v�0X��C9�~�*�cN��ۢ�����b?��F�ֆ[s��z�X\ۧj �@уѢ�ބ��ޮ�o<����������=zbTpK̵�gϙc|\bK���(�W4]�ܥ%�NȪ��.t��&h/|�����q�\���%�}�.K{�۩)�����̪H���)��ǀ��]7r;m�t'jw��\f�u�`27�u�#��_"�&W��p�.�);���P~;Wm���U=HM7�l��GLl�Hђ�����v�n?'r�U�X��6��V��}9�Fkc����j�.ښ�+{Δ�w/�}$�;�����]x�����OK��]<6�
���8Aniw�m��0���8�f3��L���N���Sj��]b��Pl�6��g�L[z��u>��n���!=eXM�x
}���ଢ�Xe{k������z��&�D���c&]�^����f����n]������@���U��c����$�*�H��7�.n�,}�ē`�Ɣ}'��� �'M��9��= b1c��ym��K�*�ۓ	kgU�໥V�j[H�
v��+4�X����Z6)&�י�B1���)�m�7�y��Ŧ�e���_�=�j��v��P��y��UȽʹ?����3��*'[�IJ�]=^ǚ<E�U���Ԉ��=Fߔ�K���\������4���o�?��U�݈�[�E\��0�_�`��jEۘ����:�M0���"���n�@�)3�y4�����]�{M��^Eg]]]�馔��>��"�8D���۷k����_c����W>���ר���p����l������Հ(��ґ�k�%�O��(�"g���tt�
�%�}�y���>���\sv����X���*�@WĹ\�\{�Kɩ�bR��*(�rwoUcMO@鴦E�:���޷c���n��d�0��W��To[�-��V�kO�m��a_F���ϰ���Z���?,#��-�� ���8�̗=_6�ٱ}���t��;���+GGl*�N%�u�\r�A���Q����ݩyyN�t��Jδ"�
$�C�W�|�1IP�׽=����-�3�_�Ҵ���]Δ�d��4!�?�$V^iRʎsK�U�sy�hS�������mQ��)??��ɜ�G�V�̬��Z����}�,
SU�!�4�t�7�\j8D'ֵ�������iZà�S�
4(���onX���X���L��{�c��׷_Z�cG����&�'SDt���oM)��TA�1�&��B�����I?N��ޚ+���N\K!RF{M�:bviP�~��b��"�W����&��Ɓ�*׾�+S�簊0!����]hh���9A>�%5��zFh�Ju�ࠣ��3H��&%޹:��(.މ9��9�((qlĦM���2V��H���週�?�]��]5��x�R����o>a����5�]u|�uZLI��A����b`�{�&x�9�zjc�MW��J�F969I��ʹƔ^����Q.�t��I���I�W��	��p(M���T�� Z���m�4S0R�M6�U��y��;4#b�T�v�g,}���?�ih�m���!�-�����m����4��v7Ŵ(���8k0hy�z�z��U�<��fl�r�N����m1D kH��4��{)����v%��\r,һj-��4��l�>����]6dG�3��&�G�ݛ%P�N%�t��)}����"@e�O�o���ܭaΰ܀:E�E4ꅻ!�����<�S+���N����d.�^����W�a��C!f-�q�Pߒ��ʑ�i������D���������Ke(6n�:u-"H��� -M٠�#.Ȍ�߃�n��"�y�w��rX�����$}�QlNV�ӯ)�&��b�9lĹ��͓�ѡ��>�nJ����Jk�%�>`�|����#�k�����0�^�7�4Gc���n�f��ף ��>n�����
r{�P�R�n���1_}{=y���l`G�&�\�4�l�e��*��	�H!pړ�3	���4f��x'<�;���m��X�S>��։(U���l(\b�7�05������.�p]�����x\�Zz�&j*�j��a�ɑE�|Ä��#e���{f^�E�YUC�׏�xq�Q.��s&Bo�����hÈ��=`��gff� x<�9�r�E&3ͣ'Q׳�X���RF�~�b�??`��8�F&��>�[���-��;o�
Z�c�m��m��m#D%itW�s�C��7�O��P0���ѓ��M�5j�8H$������(**�g���'���S���I� �#�Ine�r�/�fZb�t7<M�TUE�Q�I�1竩�[����:��XhS���YE��O����9'�4'��+bAW�~�*��T
��Sn�i�5ay�(�]�6��}��0�����hx�4��.����L�X��� �^�[�拐޽��:�����ϟ�2>*q�%��zz�b��4�ѡ�$���ܝL��S �y�,��W��N�w���ƯA����)B�>B$6��K_sI)L�ٽ��6�G���*�ga�3hQG��s�֑�.�����	�?���ҕ���}��*Q�|u�N�+��FT�B�'rt��%���b�A�ovp4.�w���6-5���V"�^���+���y\,���N��O�<*8�ǻ�'�WA�������'z���n��}R[�f�Q
~4mcG ༰��XG�U٬,/�#Ϝ(���?�`4���1/N>V���!���)����k ϳ����F��-ボ�=VH?�ѻ0CP�MS�M5���rN���<\y����\?��9j�ޅnO@�k?�2h5�RR�R��+D� �<#c�i�x�_�a�}�
��=��:;����Ι�N�r����}A�;3ӗ;���x�A%$�)��T~�'#p�`1��!��4�����H�+�m;�@EK��0��z��!-�N��E�^��~�m���eiCF�ǵA��5ǧ8���%�/���U�g�XrK����SЕ��~�����9�^��~Kv�!ں�Y똘� +N_J��`����& P[G׵8�8��+��!�/�g����.�����c��x��^;�\�.�M=�&��U��j��6�I��w��]��3>�;GG%�i".rB��?��y�?���8����������B�^�䮜���}ݩo�S"�-aD�.���xiD�u#��}�t%fj��E�w6Ǥ��vC�e�����>%S	��Q-�}��� 4���=̦�&��#E�GOo!ff���%��yd}$$�d�a�	��WSS+>�����z$��Mz۳C�Q�[��6
��>t<��r���:zT�=
~~|]]����K��#�*=�����z�^����~�,3g�5���љ��������#'-a�ϰ=4g͚�1�f���JO�RT'�uu�nmQQ�;9=mfb�l�eT|j
?ˌ�-��Zg�,��5�MѰb����������Ŷ�\���'�z(�B�=��U�\'^��a�G'4L��CJJ��h��%��4V��)#�o͕�����r��_��{|���R�j�y�M��,��=�@}���Q�_�K�آR��6sg��A~كD�*��{m�٠�_�ib�����w�PD������_�Uڵ�pp�����_o�p���;~JW��� V3̎���*���:�NLJ��q��r�=�ӿZA��?H[O�VJ`��}l�[B"T-�Q����������̬���q�-�"u`�y}}�	i�����4jH�E��9G�<�6���
�������L���D�D�ĕ��闚���m�-�y��^ȑ}��������ǹ-y6��;��}�U}������=�q�TT�����Z�1�3�=ηo�W���***��8�*�:�{݂e��,��V�19��.�����{^�̲\ke%���9���K�Z�R...%=�htrjȑ�$w}��R��sOɖ��>�cJ_������D���!�bN;Q�!���2;$|DfY�^�볻�yˊ��Q���@���}5#�����B�R�༥%ƣ��y+�dZqDī��",h~��r0�&����@ꮻ���\E�9++kؚ#/e	6�@e�g<'�;(����L^S�h�g:5��I��"�z���c�����ׯ_'$&�J��:��K�)*Q,�	/�8��K���}ww�<�[G_�c����t�<�Oٹ7�HoG���p�6�ϴ��C�K�����==y8884�/|�����<�Ҿ"��%1.|�J���HO�Wq�OB⋫�˹�S=�35-�R4����ƒ������~l�1��auu�������~�Ϥ�z�6$^��ƙPF!/%��!P<RR^�􊷲�(��� O�'�ir�O<B��|��枭�����!k��`�II2�������ZXA
r>=���1����۱ �!�fM�
޺�Kǘ��/U}yxBU�̡<C��^%�r����;l��������III�n�(����t?�E�)
���k�q	��?$��1G�(@OT�;LQC�M\^^�y��MEM�cp�sL=�J7��R����`����4;�g6f�?��ЗO<�SR*R��������/�����@u��t`��1u����.҄��%z�q[f���[W��Q����6����z�Ij�˃�Mr��q���?�a6�SD�F"Hj��2��Kv�����r��os����=����Ҳ2���ǝ$�E��HQ'�4��rzF����gWyG�S^E�Q�N#'����?V���M��І�*At���_O���z��$��HffS��|�r7xH�ʫ��0���ޫ[��WA�7,w��4�=h��jV/u��Z_͏��B��<;���זz�p!�"B��m*::�P)FJ<d�i�(��p$�Et��d\㓐��)�--+So�:���~��ax�)�5���v���,����^���V�=<Mӳ�8�	w,�����e�4�[V�HAw?���#HG������g}+)9R��.ATֈ��NН�[�i+ ��V�����mRҀ?&{�!�8H!$��qH��k+�FSW��c/�DC�(�/��Q��<�J���] ȭX�p�Xp�in�*�R���;����԰d��)L�*9n�'�#��'?�*� �Y<����,��I6���U%ϦÈ(&T�>+MX[ė@�9���Y��WNjx�t��}� �o��Q�&V���]��]((��C����ݾ�#�W�<C���_̀�.�>��BY���m�@F/��Jx��VsXT䬨������^���eŨeG�6{G�f�c�
iUmma���[�Zs�5o!zz����鉉wF�����
[������ש991���+K� �)jzec����,�1�W��N�o�+|�<@�֑�dL��&^^��)��tY<H�7�{{���3��\�9�!!!���8 HI7�)g�J����U�����`����V������:3�6�(�xqF�K��3�TUQ1FQ��6Q��迻��??���	}����VN67C,��r��A^��/|^�S�+ ����6<;3cz�Lk��5���B�"Ґ{HG���a���������ZV��×dz���rf԰����X���a�'�k�KKK��~6�{�"�����Pt��p{��X��㸊w��a;�b���4��XT� ��ZΠ�����V0�����xƢ���}CR�����`�x�U�5{�T�����n�6�I�ݢT��Zfvv5�������S-�1N�z<����0�������Y5�k��S����
�����w<;1{�w�o0�---7o<.L%iM ��2t.���ބ���x��� ��d�MTTUɣC���Cj����YY���S���XR9ق�Kj�lG��Y�M�kfE
_�R�q�QЪ<`m;����a�eͲ�ﳷ��LL�Fl}PPPM_t���}�`@W��*�����"�	��ַ�>P��/ U��B�aԀ�M��䤉���1���8���	6��a�,u�����aO��J+N6����D�<J�ڿ.[����ԁ/>�V�עƾ��?�8�� ֕X �"����y�����i ��x���l�RU- ����%�;95OV��J�?��>\�h�gVVT��Pw�m���|�̠~+GϥX���ߟ��=�ǁ��j�yr�@d�6�z�F��ّaRu^�,,R0�Mώ���t����zG��������H�+cy%��?�����P\V�lE�N���X�vEEMflYzR �E�O�tX��"i�����12r�W�`�<����V�O��]Jq�p?VW3ihi1,�=�l�R�|ka0�����f.nQy�Hp�����\��/����GB�麱�<�����@@Iep�glY�{ ���xs��mڸ��L؟(����S��Kv#e�D+���+q��wy������[�,@�,���b+���<x �ZKFN����f~�)~��R���J���ү�H+Ů��W�e�v�xui����1��.Խ��w�׷C�*��K�6�4���`����C�/� �&ef,d���,K��_���LN���;J߽Xx/�d���'�¸��s4�B�)ρI�g���J��g��(>RH�o�./�u.0Ov\�~pA�ζ������HC��/� �޼C+���q���ݥ&&&V�R�}dv�e����Fމ3�ы|�Ʉ�����-C�
�A�$�_D�[��Ha�>���,����IK��K��ɗ> ���8��xK�+���W�Z��p�		ś%��"�Me-��L燤���h��p�|��LA�8nN�ț���}����+���6&]|�8q}@�᱄� �H�~�Z���3 �_?l�G��'���q�VF�r#���fO`�F9+9�
�z��-�Ŭ����S��1J:�jcVvvv��;	���8�N��o�����Z�R�)��Sۛ(ǹ����apЎ-<*j�Y�]�o���Ʌ�+'JM���Ͼ�<g=E0�SQ��cł� �A����众<�k��R+���	����6�o��x���#	d�����s`�S=�Z��&&�{������X��a��	��׿�g����V1 ����O�z��[�����F�و�5섺�Ȃ��"X��m�b�bq�ƹ�P���������13��%Ď�L�-Y�.>Ś���6)��C��9GDD,5�i'D,����s�gga��NE�Z7J>��"����=W��t8�I��U�2���C�[)�Y�j���̆cev�`'Oâ:~�6��j`��MMHK���RPv6�Y��%�J���2j�^\�TN�˗�����o\������ �e�ms�䝕��	a��ƅ��1ܹ���w�ܜ��J3�e�xpԜl�����>�B�X��J��M�MH�37߭ �/������,�Z�%��<��lB7��K%%�Ž}k}�?)�f��FD�8y�O��77��8$�Z��({IC��^�D�H��^��>����˗/%,o��j����4��@ꤚbX�ٕ�ݜ^�Ե��F�O�.r%7�|�9��x��ͪx����ذ0��b�#�w��eHH�84�����~�BCff��/��9E��0%G��6�aa�#CDv�b�P�{Do���p�ss�Yoyv�A	!��\]/��:ҋ�G��ⱥ{HA�̩t�EC|gn>l?Q��� �XFN�^���0��&CI�TNT���E�N�xH������Z[5# 4j��V���w��Fp������q�V$��b�FF�W�pQ�������Re��˺׻���ߑL?� ��0����Ob�R �6;�T��Q���������(:R����Ng����.:Zd%wW �PMOeƣ��3G�_T��"ԸdX#lzt�q_��57{f%_��kÞ��(u�Z������t�P��˥�_wITտ��B^
QQљKǰ���~T��,+�4�H���Z=e�ީ���dsw[FKOO33��VۏT�Th�v(��Z5_��yk�[YIߏg�vjkk[�YV��*��v����+�}_�B?~����Y���[q�=%�0�C�п���IL,4HS�?��WV��v�ڶ9�����,-�٭��=�g��o��}��XL��� �������b��w/ O�$�u�4����6�����G(�I�RQ9{�fg'�8dϭ�/&�\W���>�N��#��5;���8B#`nn������L��Q�m��0ݗe�|@�������|�
���&̞���"�z�m&DA���^u�0О���cF>���V�goP��}����a������҂�@�Z��������F]r����%�;JM��=h5���`���in.a? φ'��M����	F�5o����|��*Z��К�2i\LX���NRh���|��o1))IԽc�>��0K��2�ּ����%�
z�-hA|C�T�1�&&������u qJi/t���_\�\��>�O�:�3�����
�m��[ ��*�?8\��#�q�1��k%=�3�D�"Ki�`�e.;��AXX0LݖTRz�y��E�,�!eOs]�s5 xm����g���h�����Դ��w�XS��2�2i���v�)�ZD��W�ejY�v;P�aȚ��D�������S'����
P	;īr!)1����a*�Y�3�|}���� m}I��vg��0X}m8��bv{�62:�Z���s۳㩾�{=[`�)^���R����l�{_�p}�������ӧv���F��J��#ww�W}�?�(j��'�F�m����k��N�q�왷��nὂ��ͯ��9�j�7oLML�pkEJ71�i�3��񮳜��1߿��i��l5���q}�~��+��0���1��ه���㨜���6��?�5]7�|�p����((A����1!���~��x.�
���\����Lq�����Bzp9a����D�w=�n�L̡��LpSp��o���C�Y����3�966F�7����laa����	�z�j;Hx�a�\]ծ��zZgz�<<<"ݔ
����׍�[�n����\t2�`�T���:�+ڸ��歞C>��W��Yf-�G�e�����&).�{@�ru0�x{HG����zwS����!=�d!P�O��k����ߪ��K�g�7�V �� �G4f!�*,���#)���jYE���!�ñ�5|#a��{ߔwx�IA��&���<Ѐ`I{FGVSW@<���Z�V^�YC_�3��]ǌL�-�9�dL�w�dw��mP����*nn�5OB��8>8��/; s$;��O�o|���6�!ǚy��w����9�������������
{�§7��/�ol8Ay�1�� =�-��u�|s�]|PF��n F�	X��S׶��'\��c&�/�
�9�
�E�M�8�ӷ�����EL����~�aO%�t�������ҧ?��q��'��� �]㦼sԙL�%�g�"��J�(�ư���CX duu�D�fx-0�):��:��y��T��l��#Q<�������j� A~���C!������(("_�rr�99~e�嵂J�����w����!A�V�� �a�	�����Y���B�O���J���2ܜ��P���C<I�b1�{OQ�Sx���F� '&D^N�C�Z��g{+M��%�N0�:::2=�^)aO�o\�̇d�U���į�.Bj�1�v�k����_���U���l�HS��KU������"`�$I߳���2��h����X����v ����b�˯�b�"..�q���&��r-��WWW�ޝ\"j�=��z��lP�[�l���]x�8�;���8~��QD�p���/����@���
pp<�٨�r��F�<�x�l��~��XSSS^�f�Ź "�W��N�>#%!!/y<�$S������ü�H�?�T�cb����@��q��~;�:�=�ӁW��2U\�ķ^��El�ۛ��� #z�-��ls����l����U�K���]1��v{�oE�������E!������0;���j�3sL֧j�7 ����������� ��t�T���q���I����CIq6 �w�:|#��Ͽ��Q��4lie��vŐ�/�i��f,��;�����muuu<||1�fe32YYQ�nOG�hS�JY�S�D�}	���g�WQQ�c�:n������SԁlC)�ǡ}�r ��������by�����t�U��ƃ�?KKx4��	���j��LL��J��������}����!����t(�   � �?iiA:�����n8��y���k���s�>�]{���u��Yw��c�y3'O�K�]+)���&��M�uS-�g�xE�{��n����a<b���2g˗�c07?O�U^Qa�fxǣ�Y�8����F_�A'�}��ְ(e�W�s8�b���׺�4qW'�S����8g�p���h|A	#�폾��CLN���}dt:&�!5�?���E�6'��?H^N���I�(����o�Ů��O��������q	��M������MC0I5��Yd�yb�
���r�vJ-9e�>F�	����pvO|E�!? H����eAr\��[mں,�X���������M���V �1iE(��*ɥgmU� �}��K�W0z������@)��p��B8�����n�Re��[/A9��g(n�);�;��'g��p���Ri�����ڎ���G�Z$��(51Y����^#����&4�H:�"�t&uȨE�����׽5w�Va' ����i�C��F�9��3P.��tt<���RQQ5����hڭZ'����;�wV��a�$M��|�:0���=`�ye���	����%D�oC���1c?5CZ����F����S�X�:�����1iI?~0Y��������;L�Aߩ<=�i��,��	�)V`L"��gn��vw��U44�9�o�Ian� �p�,���/,L�:W�	oUUU�r')5�H�/=c��j�f9�g��Bp0!a��O�*0��*�d0A �-/C{��!�?l澴�8A$"@��ɭ�'##�u�E�����ôؿ��M$-����W��swq���jw'�y���2qnjK33��R4"�T���W�^5��h���S������kq��ݢ�d�+v=T��_X��e��q��G*�+nd��(f5���3���~(77N����obB�D��oo�Ű3�ǌ��(r��a�E�����z�&���r�.�O@�+�48Y�9�S�>�S/.�`�5����������w���h�a��{��P�&:Pmq:�]�PS�Tد�����=���,�=�O�.#u���k麪v�4C�mݯ?�g������),,9+�N�Q�6:6V�2��&��GW�V2���)F�t���l~�"��-P��GFj�H)�牗5)����Bӄ�����^��plx8���c�H����rM��~�s`2�,j�l�w�9���g�@�i���~蛝͢!`lO8��.%F����P�u�^vc�Y�T�ggg�,��*c*�ٌ��"��X.B�
TD���
(SZ�X
m�"I=����%{�:,a���11o�÷�Z���o�4DDP�h�$''�z�(�H<��QqY���8o&��K<@S�N$�����n5j^�TRB������^�U@�F�%c?n�<c��e``���Nܑ�2��]ݔ+B���je;=}����l�����]I��(�bb��hvW7j��A�������`�����D|���)8s^ ��AY�Ԃ�#t��g�>&.F'����ØrC�ߋ��x�����`s���LJ��|����� �ה�ǃ>�;1\]]�JʍZ������P2�����G	er���|�QC*��I��L�F������ٷ�\�طo߆��`-�����v�ٸ����u���e�|[��kc��3�e#��vu0����F��@ws�ji}]tqa!��'e�I�-�
*��@�}��uj!�B�@���S�����@��uv���zt'Vy�Q�o�� ���s4����K�hWW�6�5�CDW�7��Z�]�P��_W�_�gd���C1H{��U~�����;|||]��>aN�����ۃX��DL��eq�f�H{2�i`������z%�X���ۄ�c�c������,��� �׿׵z��f��XH���62*���뛭ܪm���l�V��Ņ\(�z��3L��|���E�%����=�o�y��9͚�< ��H+��R�q�����NU��<��V�i����������Vg6P��1z�oV�Y�ە��;H�]S��p�WOW����>���M�::�#��l<<��U��j^7Ťu�p�	b��I��}n�Ui��>h"�
s���!��Va��IH���R����$;�n.|:>�@�c��.&f��(�ud#@f���dea�����R7Kv�F��RssT�-��7UL�B���v�z�]���9�<���	�B�׽���*�h@_5�����`�y�=*1QT,ՎO�@��/U�c��I'���8����/��sǓ�|�YE����w��5Z�׈�M�դ��ԣ�4s �nxP3�xS7pz<C|W>C�CVK*�/�(�F+��)�9;P�j��Z.h�Ĥ1T��uwY{q���x�]ה"�������������j����!�Ӹ�z��S���=�ؔ!�bRNM�)�{�!��8w�^T��^��]K�ح��e���R��׊���$��Q\�7�8 'Ν�zbk���i�yR#��y�Bg�����Ɔ�.����J3l����r>��r�C���[���M��Re�L�����"���կ��ܱJ?^���D^�����=%b�ؐ���(��k����Y�>�����Q�VJV�	��R[{{�A�*iu�C����["��.�W��>nN=k��j�٘!�C�I�u>�P�L�߳3��{�9�>����(e2�������r2%�'�7��ۭ`�|�oA�������Zß=9��P�st�I�O I0�i��F�.`X���p��Zl$�&a��pOF���>�!Ad���	��~�j,����X��=1;Қo�
FJPY�a�qE�����A����5tt���� �m�)��<6�£��K��$��5T�����u!�\]E?_#s�]���;�Ce��F
��a����/�V��,mlT'�R2��VD~g*�|�����1�;�ɼ3)bb�F���x_�Wo�d|'1,1�fbc�cٸ����-;[�RW<�Ou���ӓ2|��\�Gn/�N���YD0�B�b	�'�������Նģ����r?S�YilqGhVt4�e�'�s 77�T-@�����C��^wT� ˆr��᳀��eee@cW-N36�E��xj����g(z��98���q���$���4ip�Ŕ�<��'Q�X�z���}H����e��3�6�*JrH���ˆ��.��&�Ť�'���y��jcy�	��������-&5��4�; �)}�h7�#r�>I߾�o4�i���V�;;��1g��>��B�/�;�F�Y���3(��UU��h���@Ǣbc�kk ���&)��i ��Iy+46�,rVLMM���ҽ��F��:�">������H_�;��R�V5�[��y�|����C���^�����f���)=K�	�`h(���~�,�n�3?�|��V�n�*��+���q�y�8a�dw�=�k*5n�.BT�2��zǲ�y-���?]����(+����G'S��욂 Vぺ0����l����nnBUǰ�L����s��܏A���EE�+J�xxWO���B�����6s?Ш<�fU����d��K��ǎP�߼�BĢ^��D�m�vj�ZUUՖ�v�m�m�F����
����<���R�o͏��87G��� ����߀Y�z
�߾�64\A��`cg��l\���֭�@?��ȁ35��,���tJdI��+X���:������/��j���]]3�E������y=󸽽��S�~�'�}3�5��I[���單.�'OPb�iRŤ��͛=ߣ�̱����>���K�deg@��g``�,9Tfe����5sß?���n8s���>���éCJ|�1��w��3M�J�*��ܖq��U.]�BBC��,���o��X��:�geA��/5�(#&��[�Mᅕ������c�7�5��ŵ�4-.,<��^�������j�L�qq.G��LLX ��:�4���Ra���@��2y��;�[=���Tn|_w�:�G�ln��"�Y	%00P�֖ ?*:Z5BZ��ʧO�>FD@�g@r�����id��[Κ���^�AhG��Pl��i�J�������	�_��NJZ�:�an�.t�4�rGg�v��i�; ���*��R��荟]Q�ƻ�^Y�}�5�B;���qF�-�QW���SP���P\�v���IĶ��QQQ�--�`R@"Xe��A����2���hA|󙤤�uM�~õLR����%6�ӧwmmR/_���
���u��	����LU�\kGǜ�ӏ
ɏD�N6�'��ٯ�I�6�{�YRsz=��=몄BqQ57w��� �pۣ{�VHѕ�6~� ���37�t����Wn�@�N�����&���}��U�:���ٳ��{�SŃ��E{ y���+������2����{A�����C7�1H�BH!���x�~�(�1�`�5�a �C��w��לh.Ug�����2ʷ[��o�^��PƯ-���+�t�, $��b���1��NB�i�0&M�� Z�]wz*�)SQ)�Z�!���!��VQ�墾Kg�KX8$�L�D�Ǩ�s�W���QY��lh
��j�N��	���x��
�&���N��7�Y7ղ�*ԝ���3k�D���}��JJstf�������&:1��bTA�5��fffu;���\��@����JIU�gO��f$x��Z}X|�q����������EL��˭6wwvB�̴^B�d����9��3倂QQQ��iH�*����b!�ŻQ-7֋}���1���f
�?�C�RRR"

��
:e�z@�����\����aq��fMH�������6z6|���4w�E	�� P(�t]'ss�6?!�Ia�_~�.�}Ν�E�������LUU-�eT���S�w<x��-R~�0�$_���r�A��ו�w���l��Ֆ����Q�j�K3U�y�2�;O������&qps�@�(f�d��Ykt/�'��'�{";������O<%"�P�nh�aR�&�\�"m�xp�E�#nnQ�ʇ�@�nܸ�4c�7;d���Rx��E%6opO�5���U�耂奬?\I��'&��� ��*����Ţ>��,@3��J4�voS�|���p��M���W�\D�i�/��=Y1�e�q��g|��gZZT>|����7�s��$?��Wh�_�Y�Ģ���!���b�����+�YqQ�lҗtI�Ĩ��%[���=���rrs3�W�^7�φ{�QR,o�7��=U|��m����.W����Ҷ�R�ni%HA�A����%�S�=�6߬2��[}MM�{��v[/����v�P�g��X� .�}}�ł�3���@i���H<L��ʯ���]Q��e�0��!�e&H1���4[�����HߖOP�M@��U��rƖ�����f�w~NDj}xav��k^^c�Wbұ��AC�,7�rj��LݥI*Z? � �erJJ=Ո�������bc�G�|�����$��!k�&'@)�x�kX�]�l��'a�|���"r@G-=K����?	���|@�P��SL��n`"�i�����ʩ�LB���EMLLD�7h��3�*Ɉ��#񻌡׻��wBi�K�o��%̉3�n�W�QL�Ŋ&&1�yŪ����"���^�92�ٛ40����m��XM���&'u���_N��}�};�ss=�G@2��`��d���#{r������p0d�a�q�VS�lZR�ˮ����uj\�uӗ����n����̳���o"��!��V��ں����nȸo|�_G(Y�Ggc�RF5� �m�<ruz����5�O5'_�����_��#�3���g�	��EJO��^4m��7��tx�0��%6��=� r�AF��`/�vmrt�L�'X��hZ^�������ׯ�'L��J�a��B{��ٰ��<���h+�?|���5�a��#l*�}�y����bddd��$�
3���3cq����S�xdb�"k&C��]+�I3�A�xY�9���J_�m�cwZs�y0?L��y3��*(�]�@�2����񕓚���]��Q\u���ritx�W���/�PPP�a1(*����?�G�OǏK��ދ?��b�o �uo��C����GtrI��	��rS:������'Т+iG�>>��,�NN���57�P`��l��0'����׷��DI9����
�L�zzC;M���&1�2�}���'*)ٰ|��GBB���\�#�k4b��T.Degg奓��[�͟��$HHIE�ݞH���<��I.���#��VS�T��!��Vf��3���)����\�CV\u!�ݕ8ew�T��_f�Q{��\�$��G.��,�Y�%��E��8�O�~Q757��4g�14���#�轜ݏn�aa�#:�f�s��/~�PcԬֆ���fb��[e@��`y[u�t�'���PP�;;W��@�-��J��f���T�J��-��=}\���M�A`I+��uN�Y�?�r��������2.G]�����Y���4hYJ����X`^��ލ�	-�:�Ց�:�W��f�Z��0�ŘZw _l+Z���������l�\H�j���ɐ�	��Ɏ%<4�O��X��n8k�����'����(w�h�)�eCb�<��1i�f�A�����ēݞ���X�k�4��,�rϞ���Q�����V@�.o��.�镞DRh����M=�\���ٹwp0]�b��(�u�][��^��Z4v�"% ���yC���«�"���菷��ee|���C�*���P��el
T� ���9أ�:��IS�����cR��$qx��|�o߾&��=��:���t]�?�:8�&��������j�ᚗ5>{�#��t����R|�y��%Ar�K|��9u_�:�C!Y���ҧ{�����,�V���R�,YG�_�U�4��1P������ɟ;&mz(O����������J�&^c�xNM�Z�����en��q}mhNpGQ��o�)��U���Z�߸Y���X{VJ
�ĳ�R�;2l둾�3r}k�B�s�m��@G'�B�	ӻ:�H1��B�k&$H�K,�+6�+ŵ�+��-�
?����}s��� ���P�@�9��8x||}x
���R�Wvy6]ݳ��	�I��?:Ip�n�vt�D�k��[�2.�!P&���3��7[}k�.Ql�#Тs� %)	Z�C�p~~��T1�Fv�"�J/���M��?��A�jdi���NA
�C
���7��٢Kx�<i)b 6x��'_�Y+=�����������=ݕ�	oRғa�Gv���[w�\������M���@Gyҗb�v�P�3��>�Ht�,�O�|6w�Ǘr��ꛦ&	B�^b
� �����	�f�L__����t[�aruiC�@�$̤Dw山��w��~Ml��2����l_��߸�\�A>~���qs3n�ۅ+"���\gb�������Z�8]��F�"��ȿ˴���H�P*���{����r �{*T
�ŷ�@��Av��C��s�WX��\��4�����V(�+��G� ��f�_�
l�&(��T�o��zom;;�-b�]�핏��w&z�
��xTY��M��BX�}}i�Ύ���{֖@��KC�ˁ��	�,����k�
�� ��g;x�ڂ)lllx��~�������Î�||;���>�\��P_ߟC"�c�[^��k�
����____Z]U�Vz�H�b���w �?������"0����yC+��MXH�+�̤��!&�`�:99t;��$TIFFF�%*�]0H��`}+�S��PR�*'������]1�W�������28���	.N���FH���?�B}ӿ�w*K�ov$��k�ϫP���h<�ng���	�:(�1܃>�������a���k*�����AC[T4��MYYY�^Aˇ��[�M�:
x�I��*����X�S��2�ז��� X�(`���?$��u8�b��c�nZ��Տ ����wm<d��qSx�o\]]yl��rӉ�Τe;R��.;��v�������!�P�솭�;o)�	�*6�p���k\y���Gl��B���n�=攩�M��)�
���	�BQ���Rx���Z�����`��d�A��g��Sy�V��.�6��$j<���qc��$CC�T�d�脄&p�ܝwO\N��ZHI�/�@	�	.����԰��Mj���9�0u$�s��X(I�u���yI(���/�e��
��ϽֺyMKCs=R��_�4�R��M�����˚��xnvv�o��Y�7��&@�y��UWA�"�a+
怆�DTj��g ����� ÐEυ���y��������踸��z6n�t5|�N$��Q��6��汹$WSv9��e���C�PGm}o��L��%���3E;�hC������E���t K��ɴ���d5tn�`��N[8�u����kѠ���Qۈ��iH������Vl��yz�DW���+0��*I_ڠe��rr�-��x�3�gؙ�N}S@[� �<x�F�gt4 $�-���� �K�|po�x@��ҜC��V��9�˩�g�����x%��,�bQMQ�rgk�O�c���M ���A��__���M	z����@���~����z�b�"�#=��
2�r3������x��=!^����]����x����B^s(��(�]��S��-���fFF�`e�*B�_����n�|?r!tC�_����<:;;�����c��Y/��8D��jgX�h�q1h�O����%�絹���d
.Ǡl|&V����_J�1�O�n!��/�yCԂ���3빧�!�����2h*�'��$�����22�rœ0St	S���]q��!?�y�'�r�xI��Xڃ��R9�ե;���������A�(��v]� �R���N.��5,���Ə��\y��=G��CNN/��m���m�,�?����,,��K����.�M�h�f��;0��.��.zE5��c��V�;��6k���rwT)��+t� i��D���9���C�J�V�^����r�ة�	vO���d]�m^ ߳'NiG�D �??w�;r�#t��򔊌�HB~24�@&G�SQPhl�s6��������v�� E�k���c~.�o+����ZA	��u9��X�2Q��H��QnR^�W0����ѭ�g䲍s�^�~r}�^N��`
QK����+B��4��w�o_&��V�}�
��2��6��e%c���ۛ���������f�����9d�w� =����|������?��l�:_�|��龘KǓ��0�u��r���TZ�X&2\�ӛ���РJHA������:� *�NC�<�q� ����[iiiVK=ԁ[:�cX�"<�ǜPu�L��:��ώN.�#0�ƀ�6���)Eu�0���}�D @
/ꃣ�&4�K(�[𘾏v�����sn�a�����4k�����~�#�tBw�g�[K�cG��7OI�i�o����-pL���\��E�^2�F(���Dϵ�'.�!w�Mڦ�$�S򠢸���NSǽ�
	��O��f�kxק��k<��C�� 9Mi�F(�Y�|z3�TF�vUm�&�V,9Aj�*�;bbe &�{Q��>�aX�#w�J�G����?�QX������>�.�RM��,�#�6:&����=�4ş��I�Y5���ZS�8{X������ܦP�����b��3ܙc�Ȧ��?�9��������Afᕢ=\�P �u��h�s�HM����^u���"���V��l��V3��	��N���¬��n]����_�5�%�R�Z�a���?�f5ю��6���=�q%EXr�o���t{`XII��9G$�F������iǅ�q:�9'vDZ/-�V�9�բ�Y7!..B�2����H�nW;����`�0�l�>����sna����fU��Oo�����]���ezV֐��i����>]�[�����>�y��a�S��'999���������֨�D,�@���'$$g[��gff��km�JSh5]ςJy���BCC�����@i�^s�8�&�j6�$��v�\�vN N������D�ܢw>��x�����\i�Sig�/���Jb��M�_��Q�|�5�U�6�s�<��o��, �ӤLMM�y��,:�
n��Y6�����!�jx�Y4O�W�vK��=��3|'����.9?�}q� �M
�c��kc(Q��N��N�?lͱY���H��d��H��W�#�]z'�X�wd	ܔC[Q{��5��tC�oA۠���y�
j%y�[ Iӥg�\�6A�>r��#Z@���a�s�q�=p�څhy}=�ӧOF���;o���edd��U�K� ����GN��?B�Q� �9�w6[Ӱ�ۋ�up�s$��\�.}�W��s�L#_eMwZ��+X�g��[c'���W�vJ���{��!�*��E����L��U&ݛ����Kc�q�Mh���f���\�=��aee%��!��e��#������;S����]Яx~`4DD�7������������a&��\8Q��2b��[NѤ��~���Ғ��� �lV=E�I����������g�����GKSFF�f�����j�0%ep������&�`Tk�����݄�?l��������G�A�j��Qe�Z�6S��u\H	���:�a^�#�g��=���f���Lak��艉	�nkЂB �����n�:/-�F���:�H����ٍO}C�!z��YQ@֑kCy�22����p[�ͭ��P
�L8b9����=�����:��dk�`k;ֲ)_}�+MrQ�#)i��w�9ׂ����/Η6���C;�"��n��y���<��D�(��;ÙZO4ދ�ٕ�N�Y�^��E�r������o�F<��h�]���M���d��ZeZ���Q�Ҳ���(R�N&!��i�� ��u���l��̢{mng����Z]�8�|||����6���/ZZ�����m�]@������GO,�P?�()!������x�w:g�-,�A�>Th�ȬY�Ӎ���fP���w������,� ^��`����s]�]}7-��?]y���.��8Nۣ���陘���J���t�ct���321�TT�/F;������F��o� N��u5I[VQ�v�9�?ڈn/���Zp�U�&Gӑ���f%��۷{cg��|7���.�9"��[S�6`l*��$@Oj���}��x�������T��<K��[�!��-/����돊�+�W�������B4ߙ�w`�#1�=���]]]*����J�UU���uy�����N��n��<�5S`8[48�6Z"و��$�?9I5??��r�=T��Sw�sJ��8�ܠDY�}c	��N���^ǹ ֔/�B�է�꯭�k��*�de=�2!��d����rS3�����k�7^���w��sr��C�8���3�%'w��'���ޅ���V1PB�����������f�l|[��̉ʟ-�
]�`�e?iŭ*O&��5i��d+��C1�hOO�o߾�È34�gGnrO6h����K�]�蔕�ޮ�ݲ��O�y�,�0�0ҍ
*@���̓��0�^s^�ֻq㆘�>��沎�[�[K������
l�������*ÿ��\�?,t��;;;���5B#�,Zw�OU����+���t%�!a��X٥go��8�� �b�d���*�N����V������3=I����W߾}���Ls|rb����Ǐ�u���¢�n{��j�~#��5�s��ۆruD;H�k����S|����!D�5D��Rb�/)�ޤ4k���n��XX,��h���.�m5�|�_�����Z������r�f*����)�[�Ԋ���mf�2��ϟQ�L_%�݋�Ͳb��8�='��)m���lh�}3Pda5�Seg���U��/_��"����2�|\d�~
J��JJ��~١���}f<s��USR��p�;��3�5���s�<��j��q�eT��%&�������߁۳O��U�ϴ�\ܒ�ŨU2{bi��xP�sz8�\�l�p#����,���X%OW<!���������\�T�z�F�ϥ�8[u�"����r��h����0� z,��A��!g�TJ�t�S/�V��B�H��I��7���X^���2S4y�U�#�It;���e�-,,r�f&e�l�ك� �����Ykkjr<ͩЭ;�q�f��4�w�Tn<�Bŏ��/�j�>III�d(�ٯ�D�;X$���t%
S������N���+�N�R�%�R�m*�EV��⧄�w�H�b8���TASQQ�����|��maP䒂��;4�3���b�W߫�55yA	w��B����i�<�&X	;oӛ��5���T��lsJ^�
��֝��=`�A&fc��5�a�2B���L��L��L���9�c�e6��(�� ���B�W�*x���AN���aTD���###Kqs�Ngg[-DZM+mm2�� ���%K9��X�g�����}���oo��`O ߾� bN�p?9/��"ۚ��id�*j�$���D��3IԹb�@Qť��E����3���;��j����ʟ1��8�T8n������� ��Ī��M��0nְ�n����I���Z�3�3�"��2�n�y���'�U��5N�&|"���k��ђr[Ff��mg�g��2cڰ��	,"����Ї��,��U�g��%@fr^�5��ϸbX6�|��]	�K���-!$@���3�g�ZL�7�j��4HyW�44�K�26�[�o��}�Du�JW�B����ӫvvy�yl�B�*��Ku-������$�5]�;ڞwJ�=^^^��YZ^��][��p�۩i��:ԏ�D�fc��@E�{�Q֞�,))��Y�w��u�W�E���s�aa}�4���Dj�� ]i�E|���m�f�.p��B~\pӒ����(`������oYYA��4�cA۾�\5�_pd�\$�2�ݯ��r)ss�* � ��5i{$+��Q��n���Xj������'���:X%�N�22L�QɟS֨Z��8r�?��pC�/��O���&���o«W��t�D���k�Q� �1H�ٸZB�c)�[��7�M<T�aI	�߃
�f󁁭u,��Ț��V�lgg� E�b`�����u�0��)�<��'W��aB�Hg,��=;;����A��S��z��y�?�&|Hw�:�Z�8j�gc���P�'L���x\�N0���2�J��ap(a�o�l��MfFX�
9+(w@��/X����r|Oulh<ާq;��b��@�7Fk���2$�i�:��+`vTʬ�3�j�:�Ú�����[ff�.4�Dʂ�%��@�)�yp�r�����&�r�����0y�/{�sHV�WJ<y�$�.�D�����Ø�E}nmo��t@�y��A���ZDQq(w���$K,:˨͜`x/v��j�

�5��HM�+3s� ����xX�ME��,|���B�#���+[=zgmjJ;N�����7�쾵�)ȸ��偸�i��A 
9��_��)!�Am'�!σ�����ք������9�Vw�b�3;�W/%�[�a#�À������8�L��G^r�9��������jjtA��k+��k~��ۜ�_�7z^����8�:�;7J�:�_�A=`JIJ��u�����z�<	(:���F\�r����F#+p�8�q)�8�3	���.�;3G��/��AC(�:��T�.����i�o��h��n�1���z�W����A�]8<po�ꄩ���.~�XZBڋ�[7%u�XJ��b����!��jf�w���ɸ*yCNcA-|�1N�Li�O�kȏ�p�ZwH.�Fߖ���6b\ �t�\b���`�^�����P�L��I L�KL�F�r��^V�^ D�u������)����M��N�����C���L߻����ť)��CU��j7ɐD�;�3J6*tĹ���M��������u,��X\r��{���h�ZU��˝�.��9DF�H��x�<)iH]�ԁ�禍�D�[r�S�'c����b����C$/��e�����,v5�9W��Ny�Sz5�Gbk��9�y�OQ����3T�8���hs8d5g4&�)4����|�	ɏ�%2�nTt?6�h������չ���ʈ����x�����9_�Y6X���b�@���qL��=C2zXdP)��]���yv��o�x�o�7���Fx#��o�7���ƿ7�^�_�~B?R�ӓD^a�����a�	&�`�	&�`�	&����>j���WjL0�L��t���a��[R~����~b����0�L0�L0�L0�L0��oK>CEz(�G�'�����Q�ފ��נ�L0���hes�c-��R�`�	&�`�	&�`�	�?�3mF��}�������rs�n��L0�L0�L0�L0�ӿ1�j�B@<g)Dш�����p���ݻ']��� �o�&�`�	&�`�	&�`�	&�`�	&������R2�+�
L0�L0�L0��I
���X��.�`�	&��W��~AY��^&L0�L0�L0�L0�L0�{���R�wW�(���L0�L���xw����WjL0�L0�L0���1��/(c���{W�`�	&�`�	&�`�	&�`�	&�`����k#yЏ�w�W����ި��
��8��L��Z��v�L0�L0�L0�L0��/O��Kɰ����+L0�L0�L0�L�=��$D�?���&�`��ߙ�)� ��]��<����*7�P��&�`�	&�`�	&�`�	&�`�	&���z)Y�)��w�	&�`�	&������A��\�/�.�`�	&�`�	&�`�����e�W��&�`�	&�`�	&�`�	&�`�	&��=�|)YޝR������_P�>��\�/�.�`�	&�`�	&�`�	&�`�	&���z)���:��w�	&�`�	&�`�	&�`��ߔLʮ.��Z��v�L0��ѝ�{Z���Ç�x��^�e�^�Heܪ`d#&���0p�����i!�NCxO�^H�����>	&�?�Z���痡����ol�yW��W�������������������:�p�R�r��m�C�Csss���`L1��Cs�92p�G�F��g�·C�����\�"z��;76G��I��:8<���o�DGU�^�5T��L#U�	d�L;�!SLc�Q�[��#z��^�<���W���泅���c�Jt�!i�UiW�Mu�T�װ�(Ssu����n:��G�=�"�K�bˡ�ܷ��0{voc�m�k[cpe�zk�N]�ET����躹��iZ�F���VtE���՛���H}�����	Q�ȕ!u}���wln�.L�T�����:�Y&��f�\�A�mw�@����v���)��S26����'{���DI6������$��.$g�ܓk"d!ȉM�(=��⒱��pر�����+R�4��/_����7	�|��c��p���J�w?G��� �C�x�k�V��,e�K���`�����F�cZ���[�o�<L<f³���]�ŗhB�;fQA;˅���%9V�@N�eR�#Q�n��y��;S�r���{�u?t�u���H[\�I�׋T�eRH]�����}D�%��*���g`W�H�xe��\S�[��T��\��֌��l��6�=�Y�7��J5z�bi��a��{d�'<(���>σ��e������ǻ���J�E����3Ol��^[��(E,Y���ʙ��؈�L��
~�(�Ր�d�#
"O�J�T�p�YXZXq����9;��ɸ��F�u-�� �2��=�����D��3QQR�1?�B*)�D[�n6�mQ�^�s�����dC�x����jܾb�~�0�T�ˢCè{8��3������:������l@�����I���~?�j�7�p�{Jt��@gg�JX�Mi^۾���p����?�����9�芔�B��8/�Kx0\'�ݏ�mƨV��w�lV��aw,���w�UT�#��dŕ4����0ܱ�>�2?.�z�t�2;��^WSW���:{�h���J�^qT��0�Gٕ��ObZ����p���!��H:�m;�0=.(��eu�t�`H2��n~��}RV�-��X����]�Z������y?%�M����#���5�B�?%��x:��M��r�����5Q�� S�k7-؁����H���w#ׯ�&e	].�i��*��GM�r�m
qZ���o��I��>�D�߯��ש�S}���}%�._�k��\�Bف@8��q2���/&Y�⨳����M{����
s*%m�]<�E��h�z�z>��x����8�T����h����(.�ѭ+�/κ������fpHm+�msj��y-�I
�_��B�K%�d���a�;��d[���?������^��8��(��H��u֫�5�|��텕~��h�v56FZ�?X�V��ȃ~P&�	�&���|5�X��/>ݽ)�`gWd�yl�[h@���\������Yyb��h�p�aƑ?h377��r�>H9�K��@�A�"F������J��E*D[����6D�9w+��H#g~m�8�<��@6��;88����u!�bu�e��m:�D�*��R�֗�1:ܟ�_��~"�aC���$��ё�����N���0T�t��2y0����38f�)���l��#|>�ko�̗���|{Y�a*��s�l�b�e`@���'Q�Bg��A����S�F�҇wf	F�G�*!"XB.���-��_��徶[�/0��9P�#R#Q��$��-��ow:�۳��9 ��dҡ��Ч�ө�̥7�@�1p�S-!R=�������n�����L?�����zQW�*���HV�����hBv��7�$�u�D��kιv�k�NJ�'����X����ל�]�֊e �ܛ�:��Nϝ*�צ������O���hbwQh>�G}N1�m�����F�;�����5���d�z�]�[�QiQCmL�����V���q~��W�{v�2�e����-"�C��2���k~8���_���a4�(���ф��ؑ;/����st->z���<���k�fW�2������kpegg�w�4�HQ
��n�&���8�ܽ�A辬��N����&/ϴ��N=_c!��m�՟���/���x�&���<���i%Y�nn�s<��w�拇mGG�`�bC������X�޻���Y���G�ÑH�v���L�jv�d�f_�y�b�����'❶���Ú�x��Pݰ{�XR��B^���Z���č.���z����M/8=���tp�D��w�V��	�I�A:X����a�'�`��G~���"m��|?	�0˧�mf�^{�k�Η��$�L�xS��,0����^'Am���o]�M\��������g�C큛O?Tq�QJߺVD̥S��/`.�LU>SUSk�i�2��6�{=a��!�=�%����V�����{OP��y�_�����f��37��(�ڎ^>}���K�V���=�,���篤�������j*�@�RT@�4��;( @:!t���{U��K'�I��"��N@z�.��|�}���p���F`@r���k�5ל;gĕ�6�}៯�)�FA=M�|AM�9����(�77��rL��k?�������BB��t�����)���3NJ��^�7��&n}������\ɽS����d_45G�E�I�pss�]�ٹ��i�'����G�x�G�<�W��_�j]�|)�-fzx�K�8�
�{3�}hP��fl����!�/�sI����O5ǌ��=caA��?W����n�^%���f�"�����*��Bic�$����m�1��w��J���J���h�QǦ�y���w/@\�]/�Ŕ+{�v���D������=��X�s�S{����/	~��m����HJ�0���O�)G�·'S��'ml�'���!�g??�p�p�s��h��0�E@��&ja�m^��J*%����k|�� G5A
�����׹���mm{iISa}��{뒜�܅ВZ����W�e�2�Nl���$b�����;�D���J�6m(
G���V��_��kk�Q9V����㦴�����1ы�������Q�Sy���1�٧?hqKQ߄����I�;�1M�H��P�U���c=19���R� �%A=��}���l�Jː�>HK��[u�sɑ�~LR@O�}�g���ya���qީq>���� �C�OWP*�ْT��
�.�K��9�Mz:A���J� �nO��^d~����c��ӧ�A(���o������n�a�枈&��{g%�r�Z�N	۝�2�����Mӏ6�l�"C_����}�	��:q�[�.���C�G�����/����#������VϷ��2'�d��3%Eg�u��R!��Lԑ�$��͟�'�B��MG���1�� /E��_f�4�x
��4�D=L��Ώ,;8 d�[��Lv�*~��J��yyY�"��v�_3؟/al`�����%()���<*���"J�)y,ݒ}Tk��j��ZX"���u]
$���
M�I�<N�w�c�P��u����'��ʉwMEE�i�n�Fߐ�^������j)��["KP�_������GIќiE]-��b`���k���X�,Goai���򧈀@>�L���12�*�WH�T����Xj��@pۚ����gw��,�ȶ_I�34tvh��w���-z/W�FGG'�<��߇W� ��ﴜ^ijj���O$=c@�ȗ��ir	JI��eNn'v]g{x��}r1�z����|��ϯ:��W��g�SO��΍��_o,T�W�-�j�¸ZY���]���ɩP"�� ��6j��в޸���,f������V~���RRR
�bc1������;Y)�S�PH�[[��}�?"��%z�,�@)M�yv26��'��-0R�Eڣ�Ag�s�i��l_v��7)�P�Hʿ�
8��Y��O�}{T�.�5��}o��鋌� �{O�*s��?�W?X>������]�����z[�!�w�>sh.f���3,��q�=��邟)��^��iE����1ޜ�2A�Oe}�**�$�&�^t�aqDt�����^��-�cخ�޾�U��"�oM�~�zz~�#R���$	������!0=��DP�
UUUU�J��Ard���p��e�Ǟ�Յ����<�)A/MO���SQj%��N�G[�y�.�;zh�II��������+�gҔi�Z�Ҥ���<(Z�w���x��iUwww�e��0A��H�vm�������AK���i�3�D�X�޿��#��v���%g�w>J����DH(�"��@�&r(A��Υ�7h��K'�N}߾b��ڒ��H��� u�
�-��"��X����Z^��'u�����{޾�§ÊqW�s.]��\-9992(I��8$�����'xv�������Ǌ�H"d�n�9�����&_��9ބ�����Fr�b+eD�;�ܽ����6��*�q��q�Bq��'R#��*��y�o�\f���P�w_g��bL�!i�to{�)�ĳ�������њh��Cvno�u難?G�HW����2�V�cl,��4!��	�Ǐ5{b#\S��4Jpp�$�o�A�r�'W�R7�D`Y(廮������~L��VPT�Z�K˅  L����
�"������ɉ��<T���mɂu�֦�f�d�+3�1T�W��:qO��f��O�L1�esW�����e����BB�[�_���b��PT��/Sc�=��)��桫��f�~�%"b�`�����R�_Q�ȆZ�d�I[��ޞ��E.���h��u9:̷�Н�W9H���~��/!T���jJz:�����III+G� �*o�)_Kk��H���x'��;��猋>[~/�ˠ�����V��ֻ}�I�R���(=�~�n:
d��Q{�OΌb�i0��"���QV�znn�A����&(m�.F���c	3k룙��V?��io+���D�xb�`N��Td:�}�;#�%�c~{��OWޚ.o��9pN�a�6ri��x&*�Sܾŵ�C"�m������ed��Oc?���������Y,D�&���oף�8������9��.=�F[*����i&�ZU|2_<�!1�������2�x++m�6�f����]�/94��G���|�3�-�"�����r�� u2�ގ�N��������$�͟����:��p3o����ߏ�$p��wt�֓��t���%bҎ��ےP�����*(�C���*�b����8!)T@�ER����gIK���rkS)H�����������������+W�bּZ3G��z+1R���L�G�ͩ�Ϫ/]]�3�ܙ�����^�Wti),N��#F�b�X�̗���~7T�ADDDu� �gl,��?A.�;4\��;��C���������� �_�?�:C_Sϰ�#��2���| C��ڥ�����'��f �{,�BN~Ql�L��q�'�r�K�1zsz����%>ޘ�?���#x�
UdT�ې�j��I+:p+���:4Y�<�dw���(�?D�����o��ʈ��2fa�}
	�Lj�~��-�&[��?�Y�uJ���H�`{w��/�գM^��A�S��7��TLO�>=$�J�prRgg�|���ēxS�<(�`��9��c?�rH�͛��	�נWX�ĄE~\�2��}��]�=��~�|��2�r{�A$��5�JT��+�劃����r���((Vy�^Cq����u�S�Q���m�y���x����=h�	��>t�����[yI�y�/ehE�0���|�%�{��m�3��&�$�����?�J�Θ#ۖx}F/�Q7�e��ߧ�A�e�~��쭬�
���k�η��?�xL���vcs��EPg��ܗFT��¢㋁ ��A�At����PӺ�g��GOAs��Տ3�\ќ���I�5��95_wí$�`�0p�]�WE5����Z��ǯ�ə[=���㋿�Uy�����bR>T�z���۷oR�ºxq7�h�/Nw�@�(,(7���T����>?���	|MP�W���`&�g���o�����K�r�0���]y<c,Ż���^J����`�Tޏ0�>�8�C���mt]����F2��sM�[?�zBDB�%q;ȭ����(�����Q1|�ř�)#*�-s,ՠ���"���VJ�܁�~���ѝ��E��oO=�Y<��+*�#&���ƴ�N�yW��˦�{ �O"x�� ��3j�O)	���X�=�8�7�q��V�`���첀]tKi(2ƞl�Z'�x)�aަđ��s�Eu1I�J7�j�;<����:Z0��,��}%u����i�H�x�3�h.��z\@h�2Uq���r�C���Vzʰ��~�D!�znAAA�M2R�"ά���]E�V��$bY�6���ⲞVs�fIQ�=��?@b(���W`��L �+�����K,������[��v�J�������_��l������N��a(�}���R�4N��}-�݊�T\:v��녬1+a_���nF�q��z����  ��_����(a�/��.k_d����h�k/��QW@2�"ӟm7cr[�˫��Ʀ��r.F���������\!��j�V6/�"�X���Pv��D��,ȳxk{����J�D�&X��/|y��|2�Ȗv���05��o��}�<���󷶶8"8�~/;�7��N�|�^⾽�����:c=�ަ�ʄ䯸��OL���qDr]�������l�0����2�� �PI��K!z7�W2�h�N�j*ԞJ��k?~�h��%e����.T[�P<E�g׽���PN.X?���K�4��ԍ����hO@�6ƺ1���A���e�Q��\D���(����-���{1�N���s\���1��x�"+~$��y�5��Qc�B���pku��[D�����Z{'>�_~-}��ׯ�o��30�ӭX�}b�rM+P�fp�����M'���C���F���Ǟ��Jp���Wn�I5ڥ��\��D� �Nlm�j���\WP�v[�' �f�7L�b�ș�	wՁ�	#U�<9�C[5��S55u%O���l�W����F��l^�������rH�%511���	��5�ڣZ�)�:�y_fxh��f�D����&7���EW�,#0�������������7���ób��1����sJ����4�4�#��X��a�����o��QR96��kXgeM�N�H�J�x�)��xeϹ����o�qa�-� ���@�w.���������dѝ��U��s]�5}Q5ͬ�5�]�!��f�W�M�������Hy��t~������u������q3O�����fj�,F�e5����-���
��Sab"�>����q|����S�i�+;%ϸ�5+� �����l��?<�x�q�;ہf>��p3��mGp�q���6���R�#�����T��@MebT�<������{|�+k)fdם ����x�'6z�%u6��j��` �J%K�\W�k���F �&�k���9��E\?�=ʞ!�=ư��|g�X���^��|�i`T����%g�miɬ`7*�,F5]���ǘ����0�z/  �OShmm�e.��*��y�)5&%��;+��PM!ѿum Cɇ"�����{�6�c�������v҅�\|d|`
k;;�"	u��C��u	
L#�xXޗ���zu.� 6���I91��)qޞ��(#�`�[���l�9�,��"�5d����3oO���-NuqqyI����ʪK��pau�a�ꮧ��A�t�+�Rp�ոs�Kc���i�Vg?��B�&@6������X���`�HM�;?�k���k[b��;iƋ�9�3'�o�7Dr�S:rǫ��/c��~}����P����)0��/,\��j�|Y���j]�#*,^1#=c�8�"��aK,w� ���1����c >F���<�~hn� 9N��P`bJ�}��(�tf��&��1��ƭ��O�9�
�=�����ӁB��ճ�e0|[����C�v�$��vy(9�L�
G����\A�����b^�>t6��c%�&5f�9�;5y|rNNN"2~�-�\�!�\oqc�ݬ���:Cj;VŽ�O���Ĕ����0�C'>d�勼��É����!h���7�B�����X�g��|��r|f&u��5-�@K����퉘���x�u�jd�M��muI�Zl)����L�ߩ�)4��"_��ͷaz�~������p�&\���W3��������%%mK�ޕpO��@�������>W.�x�hm0Csl���]�u�?�o����{/_�lX��hx�����ˢ:��u����ُD9�o^�&��l6O�ˋ�-���%ip�C�3���ߔ2�+~��V65� ���8+���������)f���PE�� �;2���wgg?��+F*�^��gQKK����R�]C2��8� O��4ɥ���H
�s
���]�J�?[H[6hJM�v��_��(��/N|r�P��	�du����(�V�~͟��p(��Û(+��z��\��I�N�[Cl�[`7�� _�{�,�t&Ԅx�'�n~�6�Y) ��w1(��^�׳��[�f�X���E#�CW)|��eD��^�(MTDQ��U��Ѝ�E�˅���r,i���������rO��APP0b_������/��ɩe'7�7����wz��6彐6��i�b�����ꗺ�u��A�}~L�(�lC[F,u��Ս�ί���P�I�H�(�y�B��oG�s.����sM!~X���1h
�_1�<�aI�"�]���E�٘�����Qu�
��.G��F�ΰ;
���C�@5�J�x"& �X��O�8����!Z��L1��ff4�+>;Y��)�%W�4�c��/-��'CC����m���2�� `�/��U�Wn��8"�H�C?6<�t<����|vy}xy��d����r@�,P��Dh��3<̅\�0y���f������X]�|���H��Z?�"���lݪ�h�R�6/U4�$�'�1����i_X�f���	��E�׋pcu�ľ�����b�Y��:ށ� �(��~݉\���\�;��fll,�a��Suee����1i봬ɴ�kEf6�K�G�+}%�x��X��eeh%k�	{`�k�qc C�nH[���$��Dc������-q��z�T1�p!��գ�C����]�m"�^���`��L��"��}/��58׬jZ��8�Q��|�7?:2w�T^V�mq����!�XCu�t� Շ9?ɬ9�������-�B�>_-@ƃ*`I���Ӭ~~3���
MLLD��
�{*��k��s}6. ��s(?�;o"-�����L#h&�dt�/���ȇʾ���CjF�@K(��xUW��V�x+��OZ4G��\:B����Th(?�5u(2�������C����0<L�!�/N$<�&���U�q)2!���t��lq��,_BZ�oOQ��E�E��b����*�HL:� S�������A�4����Y�����4�q ungo䢚�9�xސ� ��̅Ȍ,8�*?E���F(�Λ��	�єNX���W����2���&GFF*Z}��3[�L�7�&�ߌ�����ٛ�'|���� 8��e��ȡ����B�2�����3T!5�7 �6��{{�'��W�˱��b��� ]@�r��|�_�lK]�b��eh��+*[O�� ��ۋD"5���M�������Mu"�Pqs�8��X*�1L�
ɯ��-p.����k�`c�T�j�+�ū6z��Ewc��2�_����l��w��"��I�w{}��^j�~��$�DR�vq�A4a��jv���|��d��L������#�I��9GFD����ro���3A���y�(^֒��kf�f��>~��=3�Q���Gw�ݛK]�[o�=��C��?n��J�o��~��Oo�a������V\?5���o���MU�A��q�-O��9[��*}S�05�U�������� �K��0*h�9g��1����p5��3�+�CuT�g�7Y:E����0gьC�fdq��{i��}Њ�ɽ�|~2m����L�¿ �Olk��� e��K�?V���6l����n�8�hp1��ũ~����Js�p�oB���C�Xe���X���F���钳SOMO?��Q��j��<(p�ݰ����`#�J��`������A�X��x�@���Ƈ�w��v�xݎ���޲M��<BO��{Z^�� �\��p$ZQܠ󆅅�&+�Fw
����3���`]����m(���2R�8૮u|?M��͎��q�4HR`��"{ii)�����|�G���I�Ώ�-��71�8��JV_SS��e? @��*\ �q���I�$V`Qu'��|2$��)��%\ƚ�б�yx�J3���!�]�o��c�{� � �%�DA�E.n��&��O���������9s����e?���	`{��$"��ܵ��A+�'�0��Q`x?}��/ �x04b��+.?Y�"e��a�ga	����kr��JY�f07`歭-gIVV��j���T따�����Ե��F�r"�|���,�ٽ}�T+|��>PSR��)wHG�hA��NS2����S��KJ�n�g�U!#˖׻
�x�Tq(ݻw�&#��A���S��6� $�i��>�qcY�7�;8Xz���|�2��� �P�$��i�]�o�Xı*#+��z�{��6�����ֶ����]�ّ��C	����v�ټ�>=�/�O{��uyՄ���ڎ7NSy���߹,"�!�jWDNN����|�@�,)N�U3	]��X�	iǠl�:'''+]tqKˍ�����w_�e���Q~�Y7'�d0�Ήa����q���-h������O"4]/�7��l�����AGҺg�������I����¼�=���[����Y�2�,			k8\$'v7�syxl,A\���*�xh`�H5������p��\�b�
���A�����Ʀ����"))T`����y=�jR���nt󋁯,�6oz��OQj�im�##�~z���"�W����Y(��$��-��B������s��51��VP����L���F	����(d^���<`-Z=o�k���k-��_\I�jn?cv�o�����㣭���1w8=l����6X1���N��+yR�L��Y�U0���0e`C~e�X���FW}��z|g��ѣG���$!'���j����¢���W!6I99�n����By@[��@y��k�����������h�W�Y����]���9�LS���������e�attt�Y�������6�G�t�]���Z.�����:�붏7GEݶ�������;9�0-�W5�J]�1���,�ߑ�����Q֡��"�b{{;�O(:���)^��ia�z���N8&̢
����f����+��ZZZ
k��J����>=�X�/�X�@X���^lC���I�M�2�����:P�<S��^���5�,ѕ��0�꼍��]}�8_��g�!�ƶM���WKK������uz_iF:Ǐ��ȴ��ȇ�� H$9�A￺�MD 	�m��<%�ͩ�#�vj4Z�W"M���7��fqrz�|������������C�J�\����q!~_�\l��Ӓ�+ԭ�0-��㣣�%�/?�����2ǮXz��E�%}������������/Q���~ͳ�U��\PG@�����k�� �g�$�����#'��e�>���bTT�^֡�/���,���ff����%�o�:��LC�{�R��-�n`�M�N��n�n��[�233�,�U�+:p_�&�3_��&�j�ٹ��2P���c���O���[A���(Qy�"8,	�*; 3j�֦�2�՛��#	m�c.��q��kM,.��u�,-U���E�>�a����������\�RD�4��7�?�P/*�{L�[�`�(����u���E��.+`��9�����s�O6.��V|�<߲A��iw&l��9��{ɭCS��:�	�g��ߤ���4���~Fmcn.�س%�8	�I�g��kBL0a��%ۭץ4�ov�� �NO�k���J�nc32J\�=82.ʼ�C/��{Wؙo}p{-�u��q+����_�T���y����'���Ffo���]�����c#q����z��?`�/*T����,�f�^��b]�2��B�1l񗁖[�����W�����[J�VX�2�*a�Hcn��5X� K��zh����*[s{O)i;UZJ��O��=*:��~��	AE�?&t�pA�5U�L�^Ħ�F�OW~gn�pr$��SU��oo_~6���l�{}��L�%y`��G`��T��Һ�����A
�[���"##���E�
:+E-��b̠��탍qU����MlZ��늰0��9���A��՗���S��Ƨ��::^'�a:���qbr���zw[��|&���I��5![�@�/�F����񱝭#4mL��KD+�i' U	�i�5;��~-rX��<1(���0���:i����i�>���9�,ɜ�>�x���Y&�~�|���i�S�%,+���m8r���(x&�o��v+���5ətc&}㝌�f8��0���D�#�T�H��**R;�NR9���V|&J��|?���+]۟%����K3���tbr2:�***hA�Wz̄�_WS�����J�����'B���V�r}R����L�U[�+��\�{�2bzxǫ��K��-+��ݭm6����-�詟MStUZ��,EJ\F����b�׽�9#vUMP~F?��d��fK���b�pZ���Sq��$�_i *�Я%/Ot
���\��ܒ��g}64��OF[A1�)0�~�������i�=$�3_�J
�+��_�Dn-e���вS�%僮�w����J]���ףǆ-^��8X"����.*FM߷{u�G9eeo �Cz�Cڑ0��w~|�����k����}Q�8`�Fss�7���P8f�&���:�ۦ8ݺi[P�چ��Om�6��C�X��P�ɓ��ڸQ�6��#��ݬ���7n.l��ܔ�䂷��GOe�p�:��Oe~���{@���K~n��g����\�b�����J��B��jBOJ%�&f�<8\��z*}���>�}����G��~���YԘd��r�k✜k��6�Ǜ~�NN�����~N�~�$s	q���s��,T�C�	N����='n�ſL;���D��r���+G �<-�a����?*��k�=�}$-'��#��E>������V�Y���G����lnC����J���ܵ�4�����=���������%��4�;C��&D����_Ƽ=TF�p|�e� q�岹��r�Y�g�r��|��_R7�0GUS|G~�4�A�\1�kīqm����j��^C���A�����>���G��(���İ8�+"��.'so����������j\�UUW��,=h$Cg>��f��Ը����X�r���x��v|���|$�2�qZ%qqXbXR�%���k� �m$�'n�F����}�n����n�>m��QQ���M�[�﹣�"��Kj���l�2Cͳ��Z�Q����*,���r�7��>�?ꛠy�+1�/ F��C����^�aeG�Ѽf��r�ZB���Q�m��i�;f0�ظ��\�+���Lq�OykAp�$<K�@	�1�NU:�qgW<��Zߟnwh�%ŉi���H� '����>4��i�X*�
~������}�/�,G��$�VZ�e1:7]�p9c��V���o�ϩ����m�]�:QR/+ܛG�d�=��Wjnn8���gf�����Ȃ�ֱ��oʜ۪Y|���%>��j��� F�le��)��z11���x��l�!���5��_+���PZn$�|�0	l-M��zlw��b/w��L��xN���~��� ��[��R�H<c/9��X�!���"��??s��g��	a�pj�K�C|�,5u�2�0k�V�ӄ�cGU�9Ut���j��m�� ����;����Q.��ц�7V��W�r7�\� �D�P�8ifTUM�J8�Ԡ�hu3'�|�]dо����34�w���kɖ��\o��b0���]m���p���C˓z
�G�������f<�^"	�]��$���k|��k���A��_g�H�ޗ��b�d�Pd���6̿8rr�M�0�U%�ڐ#���`\���ܢ�]�qVX������*�6y��	I5�����5P�E���<A�q\���R��*���,ۺaB0���q;�}wm� 2#JY���NS?��+���k4 }r�s�*����h�8��Tw�)�Yz�%h�3(i绦nW���Mc+j,o!/�CƤ�K �R��<9������'s�k���1M��DG"L�h]\�QX�_����3G�Z�[�s��=���F'$�� +�:U��EG��m��`���+^����v�KH���|�����  ߔS˰N!�t�1�������u����v�_��xii�w_EM
.3N���U�b� �	>�wl�	99���yz�o��Lz�iT��EM�@�t&�}��a8��Uj��Y#��%
I�\��E�ٿ���,3�;��(0���}t��Eoks�ypi�) �T����⽃�F"�Y�Byaa�c���F�n�>�}r��ip�+k����J%s.�Qɮ��]_8 �<���z��v�$/��7�u��
%ٵ��ʌ��ן!���9����
��TqGcYT=�m�i�k��?d�X�>49��f�����݉qڙ��|k������2����0zn%n�VK�4���i���2B�qI��M�ID�0+M�&�T�X�������X��jv������܅����^�����:���y�����AgU�߇��W4!0<�e��V��K�5Wll��Aϭ��"Vu2:�Χfp �)����yjZ�B��c����T2$b�茕$XkݽxaW��("*& �Qm�u7���[��;>��X3׷��.Tg���,_yzN7���uV��C��H��[��t�I��R!�����ީ?�������>��O��pq�g�#�NSYX�	o,Ui��Q��y7�B�$j�_4lr�~c���9{�~��]�%�+�6����*$�:9�<�Z��3O���ڳ��E�>a�v�����;�xtMV��D�-��$A3u��u�'\�3kc�B�������9s�tTݺ/�f̗���4�X]����le�P
$��ou�;�z����U�W�w?�(�RG"��[��П�QONl�}�򪧙��jzz( `_fx*�I�<y�ԗ����e���b1�q���lj����t�R��Cf��)����aLl>�qV��A�[s�Ĝ�;z@r?��KJf��)��#��%�h?����X	j���b��U�+��W-ς��ɸ9�猐�0��U6�Yt�Yt�֣�"&:�����g�&�@��Y�4sWHl� �A`���d2WL��,Ϫ%v�F0&&��$#!��i�ɕ�==�q
EL^�"u��ۆP��0�-	�t@�u.b3���n�<lv��P��PO�
�ҡ�cyI�\��peeD����|:ҫ� �ˬ����j^�,���4�h�cc�km1zI�R"/e�εxq'p���{�]k< DL��ȱ$�fcw���b��
����o�4�����K!g���ʫ?c�%���DM �J�5c��@�vI�sA�*�?C�O/��v�-��cd@��񿎮;>�/q���?�0��/��CJ�?�[��
������"A��9�7�7���C�ߐ�7���C�ܺ���0�i=�w'��� ���������;�G��?E�7�e�L��?PK   `��X8�Z��(  �(  /   images/52e5cf08-beef-4b5f-967f-8676d3f3880a.png�(׉PNG

   IHDR   d   K   �"�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  (�IDATx��}|�W�����WW�˒eɶ,�H���8�'N!$�&$������̓�f���ҲH�Tl���*ǖ���e��ۭo��|��˲�ya�?��~�|�93�93Gֻ>��p��Xa������^#�����X��[��ðd�z4�����Â���N�X�l�&;�Q�\ ����ڥ[pM���o-������`�{��y'Q"K3�X���V�#���+;��B���`�1C�ަo�� {��	.���E�c����D�e��v:S�6�Ug�Sð���8ÝnZOm1,�g&�%�u��{f]����ˋ��D8�+�6V  `f���<�ݎ��^����
���׆�G�QܾР��ߠ�琽�l�ȗ���^z��N STy���3c��l�Ə~�$�jԡ�~�^D�F�|�����<.�S�NYՀ�eW-�����/5lM��-]:��J4K1���u�9^Ùα*��e�ؽ�F��V�8J�3D2Rf���!	ܱ�W�ƊW���|�R�N�Q3�+��z/~�r��Q��N�@�ܗ�a�F?(�0�f�1��m}u�w�x�/pE���gՃp�v`�4g��.yn�\c��s��2�N}o�M_�7^�˵��_Ɗ�;�1��xeM*�������n�1�	�gMEm�����k2�ԗ+����X��-��̉ r�;� ����8�d�����2˝2�kR��Nk��"���0d�ZMeo�Z�ni��x<��hQp!���0�p�-�*�ܹ��#<P���Y���O�;$�1 ��ig�ak� �rm� /�˒{��Lf(}6�c��4���Z)�S�u�̈�I��k�g�O��av���O#4ԉo�&�f��#�Av1�h��j��@ԘM�j�H-�.� ���ү�hu�S_3y�ˤ���"�D��E%"{�&����l�G^�I�?Cg�����O����c}t:�ڇe�w��WpM:�_��G~W���j�/��;M'34y��,��5b���2kp16Y��F�\	���&g��1yyJ5F ny�-(�>*~�sSF�,�;�/����QX���%��s�F`T3�x3.��Kl����b�������QBΖ��v|�L�0���[n�	M-�ݍ�Y�8�W1��<x����=y�$kE�!�W�Nc4�E��s6�ܟCr�	t;"P?V{���F��ș���Ȥ�1	�ĸ�M�n��j��,�^��Pė���	�Y����k�`����Ϫ�G�ǉ3�UB_��)����gb6���-_��[��:˫l����3�]�� ��+��u�n��+��j�a��a�D�{�#֡��A1+$8�W��뇞���?IIID��49gQ����$�U� {rO��K�C��h}`*�����I�rZg�8Q���F��m�����<b�_D\�,�/l{I���ŷ�8&��l6���u��uXԛK��������s��~����1�9����k'��K���P�����0��.���8�'���v����.���v�f*��ϸ}�":��Ł�^)�C����!���<���xE���4�
�H�",P���j���X�ue",Q#3f�����*��F�YZ}ubf\� 6�_'O$��˱8�j4�֌��:�=����)���X&Y����k Q��;l�j��a���%��5-e%�*�WX�fpJR2��ٌ�Ɗ��&
���Ʋ�E�0W=��������ncs�Q�Y���!�_������"�����y^�jC$E��!���T]�9e���"�]�m��j�.]{E�N�۴���<U(�#�աT\PPz�:Ǣ,Έήf̝���B�eGB��_�����������S�����*�5��p�[������]�rQ"����ЯdB]�j8w谸�}B�>%!K��r�0k{o�#>�A�h��#xu���PQb�Z�k
���� �v���$��o��C��b�a�K��5���F���1�?_��y��P�������̨��W��~���JE{D'5��c���]���V,]�	9�/�Y.P�KrM���\���0贡�1�S{���(c��0��T�gH��)���4g'h����rx4Έ����n�j1�{Ĺ����n����X�x�2�^��w}�$.��Q^�QԪQݢX�:7�א{?�P�W<�8�zF�	��txƅ�!.��/��h����]�b��ȯ����n,xz̍솨���?뒅�=�!�B�$��ځ�H`��+�A@R����_��jn�D�[T/�\-��J�*��"���th��c߼��Z�1�[�M�����!v����}�{FMA[_4y�ީ� �D��144K�U$�Oj��rNn��m�@ThBD��ފ_4����wv,-O��E��4�j�$Gi�e��W��Ռ�D̕�%m��D!���ͬ���,/o��6JB�D�ho�O�(�ׄf_���?���g��,A��v.��T�Ѝo?}^���wbCV҄��x������*�A�"�^;d��Ć�y&k"nټ�ߍ���?�G=[����c�Q��nT՞C悥B�A�B��k},��{C�H0T��ҧC$R�0��_Gi�I�UҪU�L
�뵍j�+S�P�Hx�8�u:�v�GYޮ%�Dh���L`���dP�(��	S�g��a�����γ�{¬$l��.u�Ÿ�#����,s�ۆ�*��5`˦�bi�Cj2�I��U:l4��<����T�B�7�!�pW�C�5�!��`�I+�m������^�ώZ1�L�����.�&�Șv!~����s4Ѣ��I�ZJ։�� �;,��|���B���d��0�����+:�9���.���ߩ%�a�8�?J��{�C@hp�Jp���B�t
���4VS?��0�N ���GԽ>���3Y�	C'���cg&ʲڂ�6���	����$,@}C��yX��-"u�z!nC�����zv�.��!�~qc�&�E�B�ϥػ�����+�{�d��S�)4K���&�'�x~��k��+��,ܛ��,.d�Iܞ�6|�s�}����A!(o80aMdҤѽt�F�O.ਓ>��@ecs�H�l�<uC ��?�c�7z���!¢�fB�`�o��>^�up���}-�f�{�YM"��Tm�����,�7����}�|�|fJ�fd>�mSc������c(?BI�g�E��"���/м��N���_�Na�qq̈́���D��,�1U�oe��]�������
1�/�$F��'�V����V��B�x�f$�_ۀ^w�.�\{ϒ~^8���c 3j|_'W��#��H��B0G�L������G�x��4&_�Ͱ	a�����RT�����f2��Հ���~�X�t����9##D��
!�����&������)� �?9&����V���DEl���~���g��Z� ��)1���c�����N����g����]hҦ,��=������W��Tz�k����%�jV�Fc~��W�+_���*t�$�Ю�������1���y��iՏ"�=���߁/���m��V��s��>�R���i��کF���!�O������+5j";*}֪̍i���y�oO��|~�R�긞�6QM�Ѻ��3��ňN������엹:S�R�o����D��PQU�_D�h״�lܴ���C�s�9>����ziy%v�y��9ۼho�ǲ��8��o�%\�Ӣy,���z
�s��ݲH���4% �k)�M��;�7u�0��lM8z�ץjo�x�\���؆��!L``*�G�C��ft��m	��,���ic���cߘ���^����1"�߰p�A�#x*���@��t�͜'�$/h�\����v�՜M�:�o���jhh�o�ڦ$�g�@oo��cƨ�1*�%U�K,c�D��=�!�Q�WW�f"��-�>��+�9�h�Ck���:�x�^7y�R3�Е�b����N��
���rP����k�<�L(0k�Ȱ���|�����aD�:��M����x�%�=j�:�+�<W_4.,jz���#���ȢSV	�Fg�(z����R���	+�*�[���h8�,������%UB�9���֒������W��U��:��N��E:BƐIn�~šjM؝�ZJ���'3kX3�F�(T����=��D���(��Z�ѠӖ-_�ł�t��}���Bj���8<p���|r���wx� %���1�=���`ߋ���^,JOS��i@sSR��gę��6ek3�Ȉ/�V����żC����r�'�8|_��'r��MUC�E�����[DM�J���!ƶ�N(M�}�F0E��b~~L�5J�U)�9d��x�l"�����ۓ�Y�#,L{���љ�*�~n���^�2��"��ȯ8�fqz�3ͷv4�x��hlӋ\*jQsKX0/��bb�O����� &,��
.�"��(�]7W�+(���״[!^l�S���Xq@�O��ý�Z��<�=3Q�I�q���o��mu�7�7}^K�W7jw�Q?"3��S�]���s���z��q@�\� B��͚��EI���u���q�����z�%?�1Ô:�qq��*.*k���F�1�����ȍ4��
���y&�{���Ι]��/4e��"���u�+�����u�Eͩ'�gj��0�LL�ݫ��={����ŋ������2�?�!�@>{�1�)Ծ��菞��6�ϥ�"�����/U�y���ʑ�1a���a?�&Q<����fg�$�M�Z0�(c�k�D0�!3I7�.*�	vT ��y%9�4�����85�a��j_����w�w�b�Ix߽>&��5�j�tܭ��{ɏ��!y`K�P���+RB1��a��v���!}Ba!�b&ĪA��^=U�� F#��]�2�\|���}���j&M�S�=C-��4U�3u���Ѝ.w�z�K]���!�d�p��/k��h��y:�˕A:��ѫE'�i��0f��	z['ǋ���4�⼓L�;1'�H�°*�FTˀv�V���0y��b]}MҖd���I|��KbʤQ�0�^wD��{��Q#�kDl
�:I�����R��Rj(��r�2-^;�<g�M�	ĸ���:İ�z�q.� �_�� ��i��H����`�Ο��x���0�1e����nv"��݁��Dsw����^�fhgOl3�_�6�(Q��'����?�
J���\������_@OkД��#͂��3x�ZT7���:�=1щ~i�����Ѥ��$,9���0Q�.76۶avl8z{�ʱ����h>��[�p�������lc�=������7,8�VόjG���m��5��0�JQyIaס��Yi�R�G�H�3*���@y����b��Q`A6�\�a�6��$�QZ"b؃c�.]�ԌwWS�zT"���PTZ�7w��݁%i���?�����N踕!3�?�+������W��U7#��(�g^����ூ�/ᆆD��;/���4�i� ����P+�	�,
�~��wq��L��ߗ�����%�>�5�cXZyO�x-�*�6�O`�Xu����݊��oBqy��f�=B���xE��>��j��2B�Hٌ���&��Ivb�����*���f�^�r�d�q\�c㆕�����QVH� N�M|�������5�'��.*׭��g]C���N}M{8����ޤ:�I�q:�K&0d���j�Z�+oz�X�й:�D׫��Z��:	���Z��ܼ	Ͽ�t�P ���"v����~��œ�typX�y3�@9P6��yM�'{&�{�m6��:/��@�o�<���R�f�=0 U����~���@"3)�v�*�!X�O�vYx3��	���
^�Dq��y088�Ҳju��t�L�A��aJeY�RY�$f�x�u��fC�6(!\�`�|�Ik�R;B������Yw�>׳��FE�	��}٘�f��'"��O�����"��Њ�~]�;e�H/��t;�'�@�U?�|2�ʥړ�ę���F�%1v>��S1N�=-�f "ãq����{�l�q;X��G���/�x�6��<���z�)�Q�r9����:Q��EGļ�#R+qa�/cȞל���f�Y��gB��xf�>��^��>��k���\c���1����:_���j�=48\t��	1����bTbW�C0���'�}����V1�X���6��ڿ=SGg�bJ���J~����:���q��	�$}p�b�$lBgƖ�btV�Yztr�BprnA�^�r��Am"f�<.f��>�@�m4���B~rݞ3��gD8!\��3e�u�n�;-L����z��K�CBL~��>t����~��̸ ,2"�}�O�!J}��Gڼ��154W(G�fq�F���!��֛���mȬy��QJի�����ehܷ�na��HmG��w��Z"g�(Ӈ��@&���>�[�a&K�q�/W��u[��3���E&�j����,�c���t�~�i`at��=�VC2�[FKӀ�����As_.�+�A���U�:��]F��ybBJ)z`�I�<�2�?�)�WH+{�F�N�!S�[������X��QT*8܆��a�3�(%�Z���7�!A��4 f2h�5w� #���?6��Bf5Vu�F��r˥�V����ͬ�:;�×�`���*��b��n{t�aEZ��P:�f��H�ۃ��8�o~['9d,\�O|v�bV|L
���A�=�W�O}��j�q�V�a��kBٙR�]�U][�%31ٚ�q��ho-��
�[���#hw'�$�N��G�2�5gl���s�����X�Tܪg1�m)\|��bN��bJ��=f�:��Ix�#C_��ҏ�zb�=���D;�k��0G�>�O_���l�OK��c_������3�0��n�U�f�ݽ��O1T�!Ǡ�fH�<�{j_ŗ����,
�1��B`�u�k{=��������p�"���᝕
�y��d4�O�*�f8�`d��\q0#�E��zڊ�&�;Ž�|��0��W��C_��U3�yY\��-0<s�쯰�1#S]d^��[�S~�?�^�T�$�eI�M��sʪNa���uRǐ[��j4�V�o ��暻џ�;����i�YC��E�y�L�t������b���:�Sy�@������;��AT���z�m  `����6�jcdnH�SlN�����X4�{�1���_�v�3n,]��LGz� ^a���`�U�#��8�/t�Ԯ���N��9�J�
KK`��}v�Љ�d
cWDBL%qO֙ZJ�[)*�Q���q6�UܾD���k1�g=z����mn��E�C�Qۡ�����m�}Z�����;3���t-���w��(XPG�Ck��q�Xv}J@AnA�7D�h����v~̵~�n�����r�ۤr��hD�u!D=$��bU;�F����C�&��� �>q^���]fM �K�i�8ۙdǢ_��-5�i��O�0N�ɩ<���M[��3j���_�_��`;J뺐�~���=]�^�Uf����ݓ���ˏ#y��1W��������g>�����|��i��YN#M5E��@�x%Q�xG� ��j_%��U�n�-z,:*�6��k��{���И娶����P��U�=x`�i�=8(�nZ���lO�<�}䗕(?�y��?}7���ba�*�����_BF�#��z�j܆<tT֟�aZTyث��,���CVou�c�'�0?�[�u��3���_n2�i�TҲe�Dm0j���XF�ݩ��F`��p���O���6���A���J}Z.S,��������o��R��AN�(߇�E��7a�
Ћ���9���A�;��3�y��
��np�V�	��5��{+�l�֮Tg�=�!-	ĴP� ��|{�NR���������E�xփ���[�i[����6���~��̺E�2>�3��k���ߝ�x����)�8��M:ld�����X�3�J����9��P̜��Mhj��"��!Dl���q��\?�J˟�+T�N8c����	C��l�Boը���������W��^:��4O�-�|n� �P�k�Ƅ���:��Ħmb1Oe�.%S��K���}M&�u���gr������9����1�/�e��� �)��������)�İcb9Bo_;�SW*ߗ�9�!��!Nq�Ox�!K��kXQ^�X�N�a�&K��x�Pg�c�FD�� ����,(�Aǐ�T5q:|B�M�4��)��1'���PF$f���[�A%dI��� V���=ϞČ�}�x��Dh?�$���׾���Y�	p���Iz�~��X��5��D��L4��M3K�׬��%X��Z�}x�_��!��^��=�S�#';�)sN��ز�,�D�Ij���y��:��I"�|"+�t	a�{��П`�>1�?�|i���oL�e��?QyW�V�*&dѪ�q3�ۯ��'Mח0��,L���&S}e$i�}!�Kf$Ħ`n�b��[�U�R�T�3�?~������Z����g��F�bV^��r'�.}U��=�̆e�3㤤"w�9��ފ��
nѡ�7�X��3a豧�oލ����Db3��*�.�Җ<%��_6j�R��r]��U��1"2J�DO\Y����=q�7h�v�\Jg��^�R��Ct�;���a�FX,"��@��J�����X��v���S����Է�*[���}]���/T�����ůE��cn�u�V�֜Ņ�=|�e��������{�â��[U)@��U���+A�Q���/#���Ȟ�V�����Zq�sf�s�T���j!Ɖ&m�N��t�e����xM����8���ɭ��p����p�U��x���٢�2��'N�:��v��Twp-_��h:~y3�Q�%	�ڳK�l=�ްTU:�nߺ˸���e�O��9Ah���e�4�J^�����ɍ��y��gy�)��Dt�I�C�B���;��?�O�7�F5���w��c�b����+�"oYC1<܋����m1�^��N��ş+,�"[tSkN?mV��wU����$ﰊ9�P5�m�#L�Xt�8&PlN�ط�0����D�zվ�%��"Fbe܉�z�5��*��|7ӠEg����jtd�;.&���)��ܢ�����V�lR\*nY�)u������~�*�f�NHSu�O��M���εrl���:���a�㈊��lQh�w�;~���U^+k����Q��"����D��+��$���c�cغqn��~|�gU^,70n��V�'}�"|��Ư����z�z��~��1�3$8�]=S����	�CK*?���H��Yiظ�C�6m]u�l(��ի ���f�RrO��d#M ��-�w�%��M��ܗ��`16o�G8��|BJ�jdgnF��7���n�GO�Y='����K_X���nxހ0�IY%Nf R�E���hi��M[�����K`4�^�1��.�O��s{1�bѢ�(m�bb��7PTvr�-çj2x떭��;�9��p�n����ӯ���R�h���P�xu|���J�[����^P��K�_�uӇ�:7K��q�A��@G�HG-�ˎ"5%K�������/��)/�P�S��ՄsE�Z��/���������m���Ƶ���[{��yYJ2"��p��P�߭�3*2A$�Om�7?eBB"�At�sl��c��PP�#ؾ�'7��	y�yHΰ#���58�~�V�X�x���T��w��>���
o�������V�<���ܡ��,#��0�v2o'N�ۥ��p �n��ٮ�PO_7
Ks/.G�$�ϼ�Mu�N��)H$9a��xi�c�2o_���3t	����ǟ��ړ�������g���"2"^]38ԋs����dz^�>Ũ����Y��0�Ezٴ��m5��j���
2�7F��s�Oi�[V؏�f��+��O�����!NZ� �v
i��HW����4�x���������knR�;���Dea�!O�c�|�Uklr�Ш��|�z���g+]��u-�:�����c=���Wl�ʢ�����C-�����J��_6��<E�1    IEND�B`�PK   `��XT��"  T$  /   images/53cc934f-9b11-4097-8823-694d19808ece.png�V�W���;i�鎥YBD��n�k��NA���f���e�%�}��W�/oΙs��=sg�|�Q�@U\j\��jJ���

�(6�U����������u�N���7���]�yz[�[�x{{��9;xXZ�Z��dB��QP���+)��d�g�|��=|�͋�PT�f9+`4�P�ЋQ�[(o�>_�T�1��tj:촶�[���)���t�������O�Y���������r*����ן��j��Z��v����	����}a�JJ�,�����|~݉�ػ��qek��#��M$찮�����!�=����:���L���f\I-��i�=(����g��[I���Q'F~��6��;�c66R�M��~G<�2��}F�D%��~���ڴ6h��;�"~�f3�K�M�	����n�i�{�Ź��1�3G�A�m�b�S���L��F@̩`m���ԓhsxC�[�*���ja�b��+�" m"0��Q�M��O�x��_�f�㣹��nU�0���<���@��D���;�l�����3B�JK�P:�\=�>�{���R}<�^\�a�iiݶD�<䲡����WRl�Fյ�t�ɕ���*�7�R�b�<c�iN��L?�L�|=,u�|X���K<���5/�*�}k�S�)rߗv6�펽�E�P�kJ�v�_���h�e0o��%�H�"�ŭ��,�v���˶�z������kB��&{�+.8|6)u.^��~�rv��8p��y.(��7�z�\(�S�-z��?��T-�0Q&N<�/ٙ���i7-q�!�����{���I�Ot�2-�MLKYՈ�Ln�SI��m�ڱODsO\��3eZ$9xzeU��)㚗�,��M�pN�.$:[Z|='���3���)�����fb�ѩ���Ԣ5Wd��1�4P5�b"��Bg�!��D��A��$��'�fS�Wn?���[�+�=�����<��&?���\,���-�%&h`�W���#��9����ڄFd��>�)�ק��ݽ2��+{�a�����w����ӺS2����h��-w�̾zG� �d+���#c=�G�~�Wؾe�P�+n�����f��G=���Q��F�V�0�n>���DP#�Q.����ųN�^5i������Qc��-kA��"�����4J	Ĳ�[���k
d�I'��%W�k�k����@��b�)��H/L��rxg�CFd�S�����uEt�HEx�3D1�pU{��z]*+ޏ�Ցe����*�u%�9��	!_2)����RhY�n?��q��	46��W�Zv��T�+����i	�)5�pc�C��\ѐ8mZ#� r7{�M7������K�7繥8�I�c��n� ��:z�(f��6,tDODw����r���{��%���m����W1\��-�4k��*�"�قg�6��hp���Z0A4c�]�
E�ʩ>�8l�y�nT��S.?	���8חT_z}7
�Zs9������F�|&��焺�~�	��x�\�;���KI;Qj���Z��x�coSTM����m���H��mʂ�U֊�wn�l��]���^�"�Q��p�L��i1�*�{EX�pr�df΋u���erG�Z�k� ���A�ջ���}�pf��`���������=�h��_����	C�W<�ķ\1Nz�K�'3��U~T�0��%������u�ڀ��Oo������*���V�6O��ɂ��k3J�8�'��W	�5O�}'��^������g�$�����}���C���v�8�S	��?6����;"��C�Vn�Ba�����H��1҄�-j��%ö1���2m�D�9zˡ3�"Z1'9���-	
���v/g�J�q��`QK}hִ=�{� ��fTM���*_�0?b)�Ω�wMkO@&�ut�mf*t���늾0��d���|r6>m�AI�s6��'�-��8�����+Y��������0��a1��"�(-�͋��5����S����9 fOb5��� @����w>O?��`�~�2�0S�ؒ��1��`(L�'��K���t��?�*�K�,�ᕪDbF>�Z�F��`�y�;�A��y�tj�XXja�\l�)�b�=/�P�J��2V��56�Vk?����} �Շ�G�X��T���\��W̯k�;����ԌL^�0��ŏʥ��r��/0�Ai��@^�0���{�WM���[U\���h� s��'n<ͻ)�\Ǒ��t�b��i�H���Zf�"�9I�Q"O.�,ɗ�6���f��t�ĩUm	j߱i^���~��ïs;��������u�)�ф�]]�m��͓�4�/Ikf#�b����b��F�wk,U��D|}��>���ĔIX4�w�4���ENQ>��ShJ�MGGڸ���.��|kI� 8��0�r����qH%h�A�h)��[���)�9����F��@Ey^��k�z���^��}�_A؇!�I�i�RI�\d�(�+�#ʏk|7��V����������<P���bfG��Oĥ���L�����{<�k���^�UG|���U�y�9�����O��Ah��k���q��7�K��ܹ^�Yps��m�3x�k����#ʹ���~'���/1�yb���Mfv��9Y�����镰B�3���5�=Y|�X��C*�+�}��A/�|�\͈�%���L��n�K���~�8�A���ƨN�D�V�Ģ>�чv&�ÿ��`mjg0���?k��=,�~[_1����	:U>U�p9s^j��wa:����� �~��1��+)c.pq�Jt|lto��:�m�;�R>�hx�\�1�;��,b�y���(�*_����q�P�ﵕ^�W@��V�E���SM������5L;��ި�Y�=�ò�3�-��AwZ���L�v��A����m�D�ͳ��V�5�LV����2�\�$�{߁$�P��7���l�"��o��a� ��gfA`7L�p��K��� 6-'�7����I���)>u�����`�]��]�U�>��s�`�#02�@�;$OB��>ɩ���:]Q�t?S��<�E��N�a�UŤ��!�Ŏ����=s�I��y2e�?F�� �_�*��L��=,����;�A|C{� ��m��|^u��a�ӹ*sg��Fʼ��08�ہ�Rd<�} ����,�Ԋ�~���A`×=��ˁ闑o��2��Ϧ	�R3~r������1��{�9}�>�P����f���^	�,O��bg�ꎫL�%�X�e�k�Z0�+�xX<����7������͢�c��ĵ� �9�s"R�^BOXpWf� >�I˖����!d����O��Mr ���Н�F�&������F�D��l!�|���*t���;wZ:w��;$�e/Σ�R.D��Fl��:��st��r^M���3�q�i*C�3e��z�w6�v��,��K��g�M�
��'��]����d�j=�do!��\B�oGԴTM�߮��V��F��,�?���q̠4A��z�ƀ]֜x]���gLFFG߷��W�6�;ʪ�&�ãA�`�A7(�s{�9����f�8�uP��t�7�|��,�ĵȃH�<����w�u4�M�������\�_�i���!C�X|uyr��59�"����Q]5~���'�c;��4#�
t���o���"�4�Ee:�/t�S�|�IJ���4�G�gᵕ����1�\�ч��o�5��%�t�ة�3����'�{�
��o�˦��x�0F��|Һ��S@DQ<�^�P&����tih0�T,�����L��s�wbl,�0��Y��Z@��S��M����&I)V+\���#M�/əϮ�ɪ��6���9W��]�Hy��tnC����U�Q		L�o1G�7�,!]�Z.��$T�GO*$BLP� �$��:z��}���c�98���S8T�1,�v
$ �kn�Yh��AF���$4�͘;�;�Z��#�mUznH�^G�}�����ʀ�����[믔�G���Y��P9�|�ڙ_�m���>e:K�r��I�t����`m��a�z���>9U�~��!�W�mv˶KN��q����L� �J��:�����o�!���[���x��\�UCS�5]B^a-�p�B�ԗ���m�h��'�.�h����Q�0L�ƕI�Z��Tr���h0���ϛ�$e���7/VH��8]�
ڻ:����v�Vo}J^��/�B?�	����Y�G������L�st$�P[m�q��
y{�RYR�Njz�������K��L95n`5�sD��&���Ŏф~�ʸ���ߺ9ǻ#�b����q>.d�c�X�("�P-ç	�d�L�~B�8Gz�cή|;�ƅ�����.^��u�)m�̉9�8�k���p�^��X~z�R~z�$�_J5B�}�� bH�O7�$��~�b#�Ӱ�$>w�$�KR�|.w��=8pr�`8rX�D*@B��m�ON ���u�ܞuNb�!|��aHȑ��co@�į�+�_5�0?y��S�M���NLi��?l&k���,"�~S�u��x�2�H�C6702��J)l��]|��qO|��F��Y�@�pZ�N���|�yN�b`��>Waa��/g���0M5��	��^~k�%s�2�znf�T$�_��Tj_'�?�Y�������o5�FQ�b���C�7e��$�����~���08zǘ<'���� ׍�c?Yj�����? �4p~�>�`�>YӶG�w�$aaU�%挀&��uN��f	e�ݱ�E�Ԫ/"�߸w�B�X�̫����TX�)���4�<U`;0��=BX,�Ix�:+�s���p�%��)���Z��$����
��g�k��E�b���5��x��D�^���a�+�v�˩ax��,�&�����{J0��)U��[�R|,��I�F�.}���&�^ ���̀�\C��^�vʀ�5�R�����r��%�hU�{Z�@wpx�4��I����6&�v�p���9�K[���P'�Xm�.#kQǌ��1b������MJ,|U��O60T����F�B�g��	���H���xYPOk�p:rlE�ϕJʸ�����u������v'V�˛���r+O5�ƣ�m;��1}�$���?��Ӯ�����@s�} ̜n+�ǫ�#�]5L�g|v�©5���	E"��n��1�
��ӵ,�_����-ת��������K{g$�fI��K��e��<9�Ksa�ã��=����n�u=��|�߂I;�π�C@y���l��ʊ����N	0�t�F3�����������>d���o1������p)����|��WU�	o�f3��$xoE(�?z;�(y�#���]M�s�M������8�(��Hx���/��� �:��Y޽T���bc�c�_Rі�a��<�bad�f���9����A#5��d2�pd�Q��w�cO�_�iM���F�O�w���)R��07�b�����V�R�~�`�P&eH��r�!����*����2�?��0���l�{l5m7ȭ��V��'�ʪ��-�����s�����M���]�D�T5������V����4���;]%^�P�(��f�l��@l��e��O��ʅ�λs�����!=�Gb�i���_�0�!`.c�^rkHx�V�_��O,�qs�{u,����ጶ'3��~�{�AJ���������.+���v�������v�Z��	xKϡ�O��!@XiV��\���b��]0�BM;$���?]d��"��%�&*��Oa��f8"
#t�_�Et�#rԴ�Pp@} ���/C�㋚��fV@�.�v�':)ZXfU����MTu����2�^lm8R��o�V�ݑ�K@�i��h�5�W����[����Vp��<����䆸[���(�2�	�ר��}b�ƛ¶�cƙZ	���ڹܔ�&'^�p���L�ΖoM��p�`��6K��$�:�0J�cC^�:�6��QѷG�W��!�W�yr|ߛ��ۧE���Z�7^㘲ޝFr��S�S��.��7)�3+`�o��j�p��^�g��5�w���Ex*$�s��4?"��_��	��A���J���������ۊ،�CD����f�F6:>S	���d����#`�p�����J�2�i-ʝ�G�a�Qr����C�f7�Ol�zY+��
�}M'iN�$���P�k�:/�?l��Zq��}n� 81D�a��v��Nr����4sU���=��|�_��1����5��rcsݍ�h�1*�*l +����V�߼f�'��mLƮ��D�и�2���K0���LP5G-`�}��&�����5M'�0Wԫ��+��dm�_�GT�F㬖��OE�	��������Xel�OiDX-��妙�1��b��B!�{j��-�:��]�rƤ�Fǅ�_��/r$xتы3�9��4��'��I�8�[L�	�C��6;�#322 �H�6���������/���A�h�C9�gMI���p�F���KX�����],7R'�I�M�����;��H6��+�L��G��A����(m��+������5�)�����������h�D�˽w�G�7�n�,V�+�ktR��,����OҭD��g������}�H�lA��pf<ʂ-~X��-�^CQ����wsSn��	>����!9��"�&��h���܎���{��^����Bid���R>�EG��Ex�K�E�{��$�O��GZ��"0Wq�p}�����g�Rk!9��7h�Zߠs���ǅт�_(�}�	\��*::;:>�!dm]\TM�Ա�^<����w���<�&�Jv�ȴ��\au�:�6�ⴑ�֘�BJ�9���`��b���x�}��sۊ��A~��ĳT���9���)첊9�9��w��� ���Y#At56�d��VW<9�*�h@�B��NFQ�Zr�C��ܶ �G�`�.V�7�� �뜧���F���R����Cq�~��z~������,�>"�D;k�teW^�q|; 17�)�|��t?���P�M��EbZ��2�n=���K{��c�ƛl�<�,��FXԭ��� ���Z{��&����˲��T�;�vg7�(~�IrǛn|ߨv�|�bDC��yf��c*G�r�]���?����Kc���jcN�eM�[~�����t�pq`�Iv�]�f�����N�U�\��ЀN�.�n���6�9�5�Y�f��<*�H�@�B��T�q7�5]�/󂖏�V B�F�h�2!|d�m��G�O۰'�ޗ��GM*� HInP{Eeg �K��)��µ���XP����{��ʬ��-���/��B�E�ӛ2�F����._��+Zu;�'[ŝT_��=��g�mjQ�%#�f�e5�������Z��ˠ|�^pO������1.�7�]�#�ѿ7��~=y�[e�i�m(�p�ﵧ�w� /P��<s,$Iָ4�!�����rW�u:�P�y�_�G�=R�u�gs���$G�[����)Sn�3��%�"B_�8�� !OzWj��.�ﺞ�����ipxĚ�u��\�;�z��w�,q "7 �������(PCKnP�� �0m�Qɚn#�뭒	�#��V����g&^�Q��C�q���T}y�	��qA�LMK�~}�|�C��Ua�Ύy�jQh��?�{�)�,�ucn�I$������}��i=6p���^���:�����px'�N*"�'�Ic� �J���d�e�ʮ�����be�Y�l̞�E���Ix9�r�/r}sfm�s���3募��|v]��6P&}.au�d���X��s�j]�R����W�"���j���u���.��%�D�`��S5��>��l�D��'s����H�0�'D���;N����IpX�ʳ��1�&'�����S��.��F�pk�O��]m_N�̖.vJF�=�2��f�ga۶�f�=p)�o���W���n=��$�/����UF>�<ސ	���΁��boY!w�D�\L��輽�hqN�m�x�^w���$Mo��ִވ��|�/F[�5�%��Mww���5G��ko�cBp�KP`�|}4S=�jcU�|��"�xn�����Fz����Zh���V��&�n_�DD`��*JQ86�E�u<��0U5�>�}���tMBn�`�����L�����jQi�����P�)ؑ^��Ǯ7�.�|ܝUF��?�=6;}K�<��;�^��F*,�?�c}Kʏq�~SƝ�b/�/0(o7���ز�t4s����5Y�_)�4��'?h�P��e(N �,zp�R�j�@�?=	���$�v��vya5*o�G�M`{%���`(Ԕ��/�#yJd��5������fL��e��8�/���Ӑ�{ys��y5T㜦�#���$����rC��C���Mս� Rl�7���qd��y�O��Dk���q���=��(:-��SE��x��2��\��}����7�F�r��Y��m�4�{�I�W�!���	ggKA���=Ef k���5%5�� q�6㺁f Z@���%w���[TVZ�c$
�Hn��Z��x�T�V4�PK   `��X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   `��X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   `��X�?HU!  B#  /   images/585092fd-6de4-462f-8499-92296fb2c536.png�U�S��]:��n���	i�F�;�F:�����n���n�x����	�;s�ܹ����=s�<��@lJl   TT���� $lL��m�����EA� ���o#��hB�]R���u�~�t�0q� xxx��8ڹ��|����l�y*A	 0�+ʂ5=�N�<5g��=k�K��"3c�����s�zhj>����v8�*����U�]635����D2a���Dc������M�P~��"z3����l�Μ�ws�+<����1v��2nh���0�*�� �dz�̗.�`;7)�G�fK{�"j�R��6G��e��o���<��Z��o5І�h��+u�8oi~�'�f;- C9p�]t���F�,��0^M1��D�K��7T��*��F&���Jb��{.����a���"�P�R�9)��H��G��3qx�N��
����=��Sp�IP���=YQ#��Q-��\F�A� /R}cЩs�@} 1���H%��4�k��(6K
w�Uxt��c��[?2
��Gh 6P_�-���(�QXA1��+6o����ws��p�&E�{�Y�X��"�UPӊr�K��=1��8��K�K o��H�hV����[9�p~S��}wuZC�p=3��GPZ�d��-��jn7��~�ʸ���O�֜�����3iZ]2nT�p�'/��g�}�iU*�k�u��V��gOaG���:p�r�N�@��^\��	^������N��ś���4��Q���S��g�S4O_��&�\k����ീ�A촱4��N��u3k&lE�&K��q!� C؁HsCY��ۆ�@�[<�I����|�h5�@w��6�:<��#�w�\�ն�iI�m��G������,�}�f�ԁq�cc}�zu���'�4�6@[�KW���<��T����4.IōˍY�*��1�ف�+���R	^��>�]Ư�;W��d���tV5��C�xłyx�^hE�윽���d���7��7�S�+tP2�]��1��E�9��j����60��Aʗ}�e��3�vi#�k�cNv���� M�U����D�@E���y�̴o�U�;�]�t��n(-�"�B�}�2v?e���}�;�{��'��{�A�/7J�3�f�#��{2���t7�0����-��'@~z������
 K[���ϗYSIܯ�K�>���@ �p�^��z�k�w}�}���f�,��sT�yzU͑6�3s�7G@k��1u���ˀ�k7��q�������������>տ^���� ݔƥC��,U:V��3]�u�������&C��j!���W�>ȹ���/be\~Ii
�l+�����`$E����Χ�"����O*������|䢤W����'mo����
��glFE��_$�)�xK�EC�~H"/לiVcƁ.��4��tFNX�/��Z�3���Tlڶ��đ�Q�"F�VV��ե<_Z��������X�>��ADr�_��-��2�M��[���Y�£����R�"����R����}�$�b�E��x�@#���H>g� B�ӆ�z��F�\��@tR�>��d���9�����8������N�1~��Յ�ly�H*�n(�d5��cؑLG�s3����j=m��� 0��R�ˋT�eM�-֨�B.u&o]��?,��aGYA��i�L�s�x!�5�7�������hpy*-�l�_�FӹaQB��s��c��ٍ��4?��\�uO��`�j�!�����|*����P�嵙�1�@m�º�t�:���g(�<g�3�=��u&?�[GG �ڗ���#�ڐ4�Я)ٯ.���wޅ����0����(-�A����yC�>[}5||���[�
}	~�6T�J���9��x�x�4DE�|��_.�1�.��l�6�Gtj��;o}B��@�����̛��/R��J�q
!3�j0���[@2���}8Cv��\�MV�iM�(�L���� �G/�~S�߳����������~"���
������ߋ5�yW�O�c�2|*��[���3j.-��ބ�"���rmʅ��m����߈dd��$NQP���f�546	{���|wRZ�I)/��Pάk$�3�6����~�RfU������u�ס��R��tT�6�u��S#����zd��y�w^�Y��E�'�����H`��i�1�"+�ˍW����	��W��0r䳒s~�tC��5�n�kZ:f-��j�7��g�q����7��#M|�<����
�梕ѭ����+�E}#
�̸sૃQ�z�� Q[o�伿��:!�ޗ�qꏳL���XY��p;~��~���ΩEMBD�sw�M�!-�j8�Y��dT��k���4	����c�*[��P�4�4�.����
�o���� ����x��t��������ye�o+w��T�g��}c�;�#<�H�<geζ�����_S��R��5pVSP��{���p��7�n��P��<)�ͷH:��uj�RAҦ�(�����ݳ��/eB=�g=v�	�U���62#]75Gd��nt|l��s+��hfn�ɥ�M�N�Om�"�aTF�'?֖旱.��|H"�ǚ����ϛ�>lس�r��L���޷7	!�`US=�>4�煖W�FNú��(q�asǟ�Tc��6P����Ie���1�S"��T.���n7u!�f4����os{kW����/w*�����.��%&�b>�p%�ݾ�%ߌ���W�'����q���O�Qf�B��!n8�sn
�~j~���|7�VU�Wj;CH��99��v��\QA���o�;�S�lj�٪V��Wf4��H2�8��د38�T����ėh#�f[����M@�E�'4�Yu޹�������e��7�e�ٞ�2v�+���?=��9)��Q�#�S=Bxo�k�0֔��2��l�M'}��B�r_�f��{�7~�W����<|KD��-C�4��Uʼ�jHa�
m����ث8��N\����ZS���Vڋ��G���瞾��l��zn����'��l;�W�m�K8G	���[��?�c>H���J0�c�����;�?��w�6g��2��(�1AQ���M�y���[�d��T@�i�-����X[X�B���f�0G�k�d�_��7w���1F<�l]�>�^��M�	��q����H�KzmY�82�#�s廛��E>.&�۳�ǥ�g0c&,h���6u*����U!��2J�|^Q����9:gr�x����]-�*o�F�̱�`��E�@�Jho1N�2[�^S���Zf�:?�t���T�Řl!\X�����
�0hP�"�w{ɭ��RiDc ;a8Ir���f�[��}�o"P�'��OG&$~��4��|nj�2��oǺ��Ye��!�<?��KY�:5�+f
���ɡ�8��\����L�����/
G�C��Բ�9%vJ������X������E���7VR/A*��sBN`L�p9#�(�9���c�J 9�O����FOY��a��k�IƘ�����BpBSLI�*׷�G&��gL�a��J� .�rǥ�6�.v�_mO{拃��~_�,�a��y6��@��4m�\6���B_�	L�𣖏���g�֜疸�TüO}�>�㇁���������>��	o<ƍ�������>�x3���H��Z;�)x��t���v��h䏲�Ws��ѣM�JgBSW׻/{=�6Y�/}�G�a�|Tၸ[3��9ހD�)l��?M�7�\ա��6���]fq�;�|�0@	�/L�IZS^|�a%��Vz�����9i���G���﷞�;5o��.p����7�X`GD`t>�-�Y���0��o���h�p3��r��;z�q�����B���^�����`�vH�%�%ͭv(x��X}�c;����}`����H��yL>0�`��m���[0g��W�� )Fr�Sf�$m[Kx��z�	�۫�G%�R�O��
J��+��F�]v4�9���;I����L���8��ҍ���wN)i1j���c�T&�M"l�"��L7�7���)=\� ����z�g�a��L*t�jB�g'�:2���������2Оt�raȧR��y����8��YP�Oh���a$6�!8n����,?��C'���.�M��#����nj� �~��K�nA�;�k�u�/@G�]S(�<k�lZ��Go��Ϊ��\c�e%�d��k�1i�"�5� ��=��t?���@��ƕ�8v���wE�Y������h*����r:Ɯ?�ms����l�Rx���~���o����~�F	�cں�?�Q�U
!t�����mEE�5qs��u���2�Y���-IJ���<��&�KC�B2���ʀ�]~*IQ�%.�Q>9w+3�@^�L]���`@X4���r�Æ{2�`)��<>nLʾ�Bk0<;���yK����ޘ�J5�A����n������HƗkh�K	�%,�û��Y�K�>�b����T�֓�P� � �ΨR�V���fM�{��;/q,T ���5m��'3��6s�׼o���a�֯b-x�#��}�q�Kv�7i�O��R?@Ӣp���/'e޺"�X��ɏ�����	-�*�p%����A���
�����?��nD��@�\�f�t���7n������XϘ��h_I�ˣ�1!^hf|�VS����.�'+�?߀>��^AP�fg��w��1!蘧qs�����xAp?�Ы�㽋��`z����6�'���f:�8��l@�
˺R��l�@<*���h7�Z���<Xy�{�#���L%�v'S~W��z��T9O���gc���k�U3�@�#���U�z����WAV����S��om�:Gx����U���xEf��b�J��:��,�D���������_��a��N�(����ο^^2l����j]�������#��Z,��^t�x��&x����%�A�9W�"�{~v}����t.�����H��$�h[o_#�fá�<�,��X?hr�x�IȮPJ�n�w�����d�&�(x��L�����K��^�BQ��lc-$����mog��v��>F���}�|�S}g(n�y,�\e��C}uv�i.u�����~Rm�*��MÀ[�9Va�/��T�ę�M��0�fz�ȁ�����E<��??��3�N�+fk%�5z
?�#f�(�*�����z��'�EH�
�:pơ���3tL-�?� ףg�Y	�h�wq3�wY��Ë�R\�d�{�����c{|���㄂<����/S��Y���f������,��C_�Y���Sm���ay��.cy`�n�͘����!Z*L݌����63�us3ˣ�c ��ݵ�h�~C%�A-�.�&��`Ƀi�U�H�*�~r,��i�'a����ӂ�����k,eFJ�`w�5o+���D|d�ɰ�KP��d�:M�`q��~���H�@K�y��@� �cidf�_�=c��`�b�yJ��-O�8k}��b}x@���Qr�bIi�\P3��,�a�!�_s�����K<����v�y;��j�WU�4 {��}N�b��&�$dL8�[c
������*�ܙ�8�B#F4�F$��*�~ᚾ>�IL��D\��7�6y�lHY�E��C)3%�᝶�nzl��ë&�G�$&Փ�B���'�`l *#��͙G��i�7dij�ߟ36�Fs��e
��xW�<Jj�i�y��꣰`\�H��b$����;�c�V��DRŷ	��\U��ͭ��y�آÚ,x�{��K��R?��E %�GU���:i�@Z�H�������٥�o�r������p��9m84!��9��q�P;���c������q�N���`�<�_m�_-�O�}�w\�N�Z6���ƾ�M��՞�������Dٙ�b/�BW�M�XT�8�y�����8CKі���8�h���T/\T
O�Z�V�L=��x���,��x�v����J%D�����i��[]^,��G�����>z�I1�E����'[�4kq����((fܒk�x�`�9�Ń�7⏑�Z/t1�$W���{�t��s���ܠ�UO�s"i���'�X3���>2�������O��j�#�]!���IhJ�D<]���������I�81��2��6�|q�iǂ<���Nr��;9w�=������8,�X�&p`	��9w\
VG.�8.q�EM�iY���@��q�1m�j߅6�}�	��Q��su��`�w�Q�i�[�l�!fg�>��m���wM$D^��+|>:��˖ޫ��Yߝ.6K�=0č�ө��e���h�s�{���x\��Y���*�f����\r.�
DQy:���[t(5�jM���d$���K� l#5�wǐ!��ɿ��Y��D*��;!��!9�wŲ)��
]�Q	�ֿ�/��q���������!H6���U�o>1��A*CP|�g����)v�J�������~A.-�rE�6.�(����$.���H�)�#t�U��+� �G����_��?���/�~��fO��)|rn~���S�Fo�7���R5��|���:�?N�d��b���g*-J�[�'ʺΝ�V���0��KӠ��K&H�'�������V����!��rC����ڳ˸��|5i�r$KȳA$��r�h�P�-T�'z�g��@�H`�;�<)�E�>��%^�H�6����n�����M���r�\�h}�*��V�4��Q�	����G������AR�M��G!N����v/0�����zy�����Q�!�WNqY
��o�04m�[�9�qQp��o�W�fSB(Ku��#�<'��'ϭ��gB�_0pA�bٝݪW�FX�l��I��N���2�&�?�����0(�P����=]D[�>302lv��̫��<⍌�^¤��q�Z�О���Jі�H�⿷~��[>�U�R lļ�R$y��!*�(ǻa@}Ne��`&<�!�I�ʐ���ć��m����+�&@�E'Hz9b�o&�R���&-�v�hyA��<�}B���Ҥg�(�!�%�jCP!G�jNnnD���ژd���.Π�i�U7L����\[���	.����!�A�{ Q�Y��?m��ak��f�1.00�S��!�sSA��f�%�Np��(�����-<��t�d ��0���	j�$L;j��
�\�p���ڱ�������{#8�x�ˌjN�TnU��f4��u�o�9�uD����F<R��e~�>�Kb���$3���D��x�漹��h��x4��a@������_Fc-�(��7���O h?��~I+6�~��/���h�Y�i��_�A	�������eT�$Ўl�U�3:
U:�P��W�6=��8K�V��7yѰ�*��$C�O�d�J�D-��M�S>EKN�*%Y9*�B絥���*7'n�JI`�CFʄ�w�����	C�:�.WP��1%�3	�[�lC�V��G�;�h�Pd��]4G���P��l4�=@��2����?�#N��µ��F��!_�Sm�4����dY���+w��V�r;�Ovd=X�~ɠd�3(,�WtL�jG|��/�B>�Gi}%聖3�1�T`~�#$���I��a��AN�'���,|bHM�3�-�"_�_4��1|���P��8E����,�@J��X*[)<߁�2���r��B�¼#�a�=�%ە��A�Wߝݷ8�^F7�fz��R�b�M�n-�k�A��\t��_P՜~f�MG'�sg������Rn�7�Ѻ����"��6�5�;(���~A�nԹ�
���s��6ݑ�����Z&� ���c�I�y�?�l����ђA$�͟��9ȧ���f��cPUg��	(u�>#
㏾��	gA̡ɁX΄ZcX.砮���hT~Q�v�z#���ph��'7��Z��Y��Z"��Y���b��p��2�s����hS5/W���G�h
=�=ZY5'���4��3�����WY'�����,Cf����d�:���*���#�W%��W�x�s��_U�I�홗�����1\)�e�Er,s5�r��YH�H�q�1û��@2D�R6���
�6y`jWDA2+9���Kf�L��9l.LU��v.�@�����x����X��񪼗c��`2�(	�N/΁����΃B�,��F9S8m[����Jq[�07w,+��
zE>�M@}����V� K�ZspK�	�щ����M݈�D�-MiuQ�|g�9{ٝ��|�C�o�k�n��Xdy*@��*m�����R�g�1R-Ks���9�d��j=s1�m��x�sms�O�1��[��Te+!�A�PK   `��X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   `��X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   `��XXs�銙 � /   images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngl�T�m�6<Cw�t�Hݠ�(�(�H�H�HK�tww*#Hw)=4���>�s�k��Z,��c�s���M���2>5  �WUQ� З  �\,�'�~��oh.r�����/�E8�gl' �������.�C*WE}W]GKW����l]>�;}�u�l��� �
��=3�=<���1���/�U�Qq��hZ���DĊ2d��s>�u>EYẼ�SP����L�H:���pt� ;�y�o���P(C ���ȁ��e�$���)Й%vݚ �������f< �٭�=���:*�������0J��	���� Ԙ *@F��u��}$�)IzFf�Y�	��$��;��8d�+9������%F��-լ�u���{إk�o]s���W[�Zx��d�Y�9��$����ʹ��R����a�%燷[�2S������x�9�w;2z6,���2���� H���m�z�#�2"(���	�X�w� �/�q�լi<hk��.��\�X��$O�߉��s�g(�4'eh�j�w����Pښ�ᣔ��'�K�sI�NY7?ι�X^��2����D����/�<2��|�|���F��i�ŅƮ����5�H�Y+u�7	з\��NC�/�����dJ���:�^� z71���'"��gl�n$�n;{��h�t����u��va�"��bEie*�S�c�#m�t${F�滬�k�уQ�9��v��@�MW&~�[��l��Kl7��v�^ݧC�>-x5����n���,��XQ,�����Od:/z�γ��Z���Ol[��k�c�,.&�� �U��"���mކW�L�x0
�����w���MZ��P�0��-R) U2o�Ng�����dt40�R�r<�:��qݦ��L�,%]�+�ä��SvxA�mc��}��O�C�Φ�U�$�b>3�\t4 (gn���'`{�'7|�K��h
`h�F��[Q$*��4����@����d���55�y���=��$��n��NmgD�85f����!oc���_ز� 9L��)�)��1��G������ڈ�x�N��m�0e��/�-Ħ��T1ɝ˟p^"���� ²hHF.>M�<�n��C�#�d��YT������sۅSV�Zx�������fwD�ԼX�n������4z9���|�����e�2�hC�~L��c��Z�¢}�Ο�7o%�ð绡�p��}�v�=3�M���� v3o@�R��:�i�'^"������e)��u�����_�J2��R�d8��'�s:*�U[kj���_h>��gr����͛<K�>sN1	H�=0Y�r���{����$�^e`�E��"d4,�S	?��� x>{�_;�˚ě��������X�J��T2A�@�'�K�P$��Y���e�R�l�MR�$R�㺪B= ���o��EZ��8K��`�$�40���Cˊ@1\�Y�ӿ���'��-��e�Y{����Cv�:�m�V��o����mj��Ԑh>qz�'!j(�KO����gn4��JyC3�M��?��"��`��M}\����{�\{t\S.j�3Sst�߫��/�8T���3G����6�gj6����O�0�=�EЏP�A�v�#I�����>�����e�|��}�N	��¿���#��+ ��RY������/��W���K��\,����u�>�u�mUx�N��&�n���K�*ޙ{�L�e]]�˹���M���Jюt�+��^<y_e�<�[2{�8����@��AbZ�k٠<�:��V\����A������/�5EGg1c}	��=���%��~�ߍR��p�f/i~"�T�>�O��:�� tw��f�A/9�۽�d3K�X����mh
���_aߒ���;��^��˻1$~ZJ���}�rz�=p�e��w��/q��)�G��ބ��[�u��](�l��g��w^�8���tA��I
je���R,.t#�o�b+��ڔ�7����u��H<�I'�g�����(��Z~Nv�5��h]�1F�R�Ç�pw�$sC�6$K��q������t�ܭ��:Uq�-�AQ����?Ni5E��|�o�ڭ�5 �Ǩɿ睳���3ﵠ��� �ݓ��Aj�s�>��t�v;��\�����;�d��J֮�����P�8�-�{���Yz�OMGi��Z�������O�'�{�Ute�P@b��fO�C̷y�8c@���:�������M�G�X���6dտk\E�j����l�dʛʴ�/e@��0����o��8N��
���]x�)���5���!p~�i����-3���Р/8�r����>}m�#�4�1��A܍	;�0�-�M��a���%�� G�<����6��`ȏ5مt��u�WtF��{vhb�Ѝ10�h��	��A0� F,����4r�@;�Z��"ŎI�]�[e6�ޟ.�.�v�v����x}R<�_�)2���Ǒ~���ms!"�(>p��:g;������(��E�n*�����c�ͽ�k�mD���3Z��&��s^���p�e��d^�36,�sl[��S�8��U�+��_����EC������?r�٫�3�Lf��,m41��[��@��a��偳�/T�N���H0�F��v�6��8_�)"c�J+H�ǋ�;�u��@XƣF���������������i��$�ͧ.�<E��FbH��Y�t#�I��C����XJ�Ya�a60��p�:��޾�B���Ft�G�\��~_q��4�~�_Y�rt�/�D�8$��Y&d(�e��)z�po�sqA���/w"���/,�ܝrWC[X|8�����9p�LT�������O��7_�8��vd7�����~zN��+���E!�V�F��_���r��m�m{_&�z����˄�F�7;��+t��i��K��
�>`Xei^K������'N�Yh�W�D�&"��ٌ��yQ4%� �G$�K�?�yw}G9h	d1e�����-�<�:n0�x�;?���@������\ڶ�~B���l7���[A��ޫ'��g��љU~�B��㭊Ac~x����z���,ɼ	D�%m��廓��j"�x;X��|��4������]q�{fY'��;�,h��fe{�[��(!����L�b�=EϬ��δȏ��۫G@�Ԙ4�KJ=�9n<ߵ���hu\��uG;�d�/]�-�)W��NqB�E����d�]Ha#�?J��c�F��zZ ?�]���c,���VL"zlO�1*�&~mMݫK9Qw����S�K뎿�_I~r�g�c���m��)z��D�6֝������M�b�0���.�q�5�ܑ_��O5�>𩫅�'o"kE�]�q|�u׾����s��"3Wz���Dv�#N��G&qz/څ�U���P -+�k#���7=���Omݚ���%X�m̭��`�f[��̋�X�#|�!�������j�H:�j� ���$��9���2����l�8�#{VQ���$����I�Id:ȊI�.��)�����?����d30Naպ� �C�
���;:p,��׫�$`�13������SL��׈�j��[�Ƶ���wz���y/~X,�2v%Ae�[s�=�Bs�ܦQ�7�f�v�w�
���p=ח�N$b��+`ǹ��B2�;�،�ƛᲱ2S⋢����S�[�%���T�d����0�װo����>��}�b�w�t���4��F��kw��@�Ad�}�<��cmΖ�seʈ��O�w�\ľn����%eR��KLli� �5�C0	k5L�����I� �����A��i,茽YS|<�,L����e�hX��Tx�.�Rqd:��ғ��t��4�E����K
���ʀ���
b����AF.v��FV� ��Ewz}j�i��T�sz2Q��,c�QEY�e������lG�E}%���Oz� ��!���$_C���Q���ǃ�O��r?����1��6��W����u؇��L�����;u��zco69\h=���1)��}}�!�\׺m�28s�fVes����RNb+��>R����U�ǉ��'�4~ :*	*ޚ�+gϥ���S~v�$��-�Z?��O^�{�,��B]��@JC�����(�:�ެ�/V4-~�`I��9��c��
���ײ����X�k@� �m��q{&]�
�����Lp��_�KJ8�9�)tc�Ke�ےϔkl� �w&���d�UZ��I|��)H0Q��A��Zry>���ˊ˽�y1H���|�T�g�<����[�Xe�>mC���~�~ؕ��sz�������E+56Џ#\���L�X�>��d���o���/����E@Q��Wid�-� qt�n�y��+����X.mԚ��yҲ�d��l��B���]S"�&? }�䑑�M�޵�^��ؖwU�e,���h>b�?\�!���Ҍ��e���N1mqz^b�J��.��+D'j��(����n�(�O�[��;W�}����r��А�+����U��xI����������Q��9��[_�[�x����RUi���./��^��N��1=��~��;(݅Y�:Etl���(���� �̠1 �|$<80$K]j�ݰ6|`��x��L�)	o�td�<��P�{5OA�g��ݜ��72�,>�H�2Gz�x��k�2C+�/7�`��|�^p�fvڕ�l�3bVr���<]m�ø�W� ~GNV��z�#���"��LΜZ����1&gI��O���L~�j[��c.�e?�
��kMS��G�)�<e6နO�V�W���C�D��qL��E���ic��䯗����{�n>������˕H?�
��	�/�	�̽���3�i���:8{<��B[m9���=&YI�,�B��iz��<�=	���X�l����� �	�f8��1Dߔ�zޥ8M��T͔��tߤ������Kk�o��i��䳸���r���l?`� �5|��G�y#���*�i>ɒ�?}�'�N���2���֙���I����γ�兛dmB���ӟ�c��f-�<����'�[d�fzX��|B�����ϙw5�@v�c�~u�z�c��L�F�~�rd2\���d}��"�����9:}�I/w���)���L� �0@5c���z�.yϟ�c3od�N嫮��u�d=d6�囗��a�v����!�w�ܞ�)1s�u1�2�Ѥ��@�id�T�6�%i�Ef���ﴞ�U_d�k.��>Q$rz���gؽ��S�SQ���u��>��.6��1WvsKnsK9!��dZ�_��/e��$�wC�|��
�(��y�f�e9ܲ.:��l[�V��~�㸄V�IH�vvn��[~�/S���jyСl �jf��y�2>(�=�����&H\��%���{��t��	=�8��G֝�WP0?����/ ���o����d����ߋ9��\:��7�c�H^6x@�!;[?���v|�RC��1��R�& k�S�ud/�'3m����($U�L�'�Yh�����lCx�xƛ�֐���Q&\��U��TG�!-�5i���X��O��o<�B�u-�%�O:�C(�S��v�"{���͗���B݃W��W�)��?{���!��u5���>��7��dG]�r)b!+�AQ��>3q��VO����2!cPϕFv2�즪Ө(p���ӂ;v��/���S+�����J��?�0�Qj�u��xF�Q�R�c����HA:|�u�J�u����'Qe��7Ue�;"D�nL�f~4�M�5�1��l���2CX0��ݰb����E_�l��9��L��A˰��k�� �Ar����uzG�ӳ5��aQ 2��/t�j��5p�LF�i��YD�;�N
 �5chŏ�x>G'�hQ�9�L��uK�u���&���Y�t��[�f,J�M|�X��S�)9�;߄ĦD���C�Ԡ����a��y[�%��v���*�p)W�D�f�Q���a.XM4ף���{D�O@"V���Q;���������}��^��ɪO��hf)�gG��_��Nۋ�%��+��Tq�;?�c��'.��т~-��W��T�05)OpYփt�
L^��\�\mw�@���'k�Y���8�߄�Ғpy��A�R��*G�|M�h`�,�l5<����	�	h��/�Kr��"��A'�W������x���$N^,��0���؝�i����Xr�w=���*���Or[s��{�>;tI���E0��?�7��9j�R�p�)O=�f�U^�B&,��D°]w���O�tz�/�AoE�=<��d�%������+�Zд4����~�Q;I��
"�DM,�����أf������p�U�+�/\�L�^q���eGY���N��/qh�cKHwmC2%']�L�:0�Fe��f9��	 �&t���0o	�����)tZ�4�K�]�<���K�t���	c���߬�3F��K�(�<��%�bՖ�#J�齷%�@*���>�� ��#$�􆼝��&%���1���)&i��Z��`+w5��:ݍ���*f��ѿ�d�|?3,Ji�b���<^T����p�ņk��0�|����ۡ��܋S�W�>}>�y��+���v�#Ba�h�0��,�0�q��)�[�l���Dis$�)$>��7|�o*�X���?|9Gf?W]�ovmmJ��'ZW�HJ�bC�xٶ��\ \cNU<t�L���Z:ª���+��6k���v	�j�[����� K*5�`���	h�U7��S��]���1�o /���6kf��U9�J�;��Ӣ� o��`�>���4Ma�hd�`�_���2���\�Z�����ϸ���*^�]?lӎ��$�-�h��R�u�H�r����� ������bv�?�WU-�nV���d���w�T5�\JH���]XL徂����('��5ֈ�z���jjK�Y����Cr�����V1�rE����|)mR��4�m!	W����j{Z Bui(5w��lg���5뺂V~����8���k����#�ꜻUGe�U ��=}���+�U��q�`l��)��k���r�g4�ŕ��M��N�����5�E�1-�	%H0���'��Ƴ�A�{�9�C�����nf�,���cm2U��yI���c
.�T������7��F��R��3�u˪�d�h��ڋ�υ%Ju��}$S���D�	�&���,286X�5#G�q�>4)?{Q��.�ۋЎ8
�	>����:�] �̬�q�owZ�:�u��-�m݈8��� ������D�ñ��Ñz]i��l�"�[��?������k$��S׾���:�k"�
��w����& 	"T��
��۔�$T�h4/15�Z�Q���Fl�K��!An��ݷP~6���TPp�E9�W[ـVT�F��'|(��n��3ռL�e��}��짢�Ds��SK&��m��(�	t�j:ۦ"��.�m��aU�x�d�\��^.�����_�w�ӓ�dS�g/Cj`���_LB�:�m�F3�pd�M�C�����i��o>�Db��J��d�+B4N
��]&�;�ߠ�1C������z��.���l*3\���'8h�Ǒ)A���l)T��E0mT�᳑���;e���5:����N껫Wo�Yr}�����s9\6�>dj�T�xfd��^�=9��;��[��x��ONQ���E�3i�k�x�9�l���[e��O�4hl�e�_�QST�҄�����+�"�2n�j�F᎑�$��T��j���e�Q�"�H��wl����~so ���+����4׏�:���ʦ+�缬2k� d�M Bm�,�ΦMq��a��W��}B���BkM�;����;x��B_�㻢�>u��D�7�������ז�`Rk�H-)R��y�#N��	;sUFt�ө�6�$��Ƙ(X�葚�@����[����Y$m��Z�oK9?^�lgdOk� ǂ�
7?2StF4�[���n�pv����Ҷa�с�y�q#R+�)6�t+k>x�ѧ��ϰ�zQ���h8�55�sf1Qvk�v8�K�D�%�%!�.�G���|�HO,'����o��k�1��Ntdj�c�2@QY��S���^d��5�AH���a)W:/3�������P����=D����PK�G��CF��J�yk.��f��a�N�>�<H��(�z��8�!��M��vD���4Ř�Q6��Ӹ�	 (ԏ�Ea���������s	��"Ζ����!9N�q���)@���T����l]��i�;����u׹�K����ƺ]�>��7���e��^6�,ҷm]{
w��(�[���J2`���A>,����-%Rd}��.�G����QSP�R\�Ʀ}��E���y�)��)�ζ����֩����D~vO�[G�m7���<���a���H1���������q��������佌0�rdP�`m����c�e�O-����b��:�x�o]��C��ĻDs�$\Z+T��ij��;J=#F(����+%�(Mtej����o�U���e���"�%6q�C�F��q�L�__ѳ�y,[�o C~b�O��b��q��5̤��B���1:ZU�����|Ij�1&��xlj樝f��y\k��Ñ$�ʄ$��XQA}���گh��3��_����D��!h{h�zYO��l_����9P��m\�R0�F�y@�.!_.�k=]j��>8%�%�,]Ğ� ���+/Σ���̜�5����r��uL��r ��7Sc��:��0~T�p,L4�r�еSW�b�S�=#���Mô-��D�}�eؽy{@in����F������|��W��@TG�j�ͭ�9}܉���q�<�8����`�?X~-�q��U����%�D�39+�x��Rb��-^�:>�������;
"PყK!˻ER�5M)�r���l<�YD��w����p݁OZ).��A���S��s�D�Ɋ��ЁK!�␍*O-���s�{Ƚ����w�s0�s�kB�!&pfh����I'A%�1Z2�Or�\�]��j4�j�������-y%�%�o�K�b�H�}7\,��7����̡�M*F8������>�fM	y3]��'�zry9ǎ��sP���ђ�#�<��A���J�N��'Th����Wna������s���jѽ������9�))����l6�/!�m2D�mM��f�%F�d�#�O��ZoE�WQ;q\BP���u�t���)����l�z�7�ެ�)/-�s� �^�hH �����6�h�W�\Tյ~HS6��Y�ktl)��1l�z�������I�E�h~�5���殜;�;����i�衴3;�r�`υa�1 ��R���$A�[�%e}�fMQ)՝���hǉ۽��t��B���[�t�x/��
�����u�y��d� XU�n���H��S_,>jۥ|�?>@/������խg`�F�8�dy�2���_�bd��Q*2�xn:ۢ�d:���|�ޥ��L|��R1C9���9���;B}�l-.0�y������q�/d#�ц���4��o0���Tr��'B�����~2Nt�=1�[�a�Ù�bCx�[,>�M�lٱA67���,���oxĞ/����Db}��}�;����,}=u�_Q<`��|h���?����^r�3'���'����W��d#��o��
�}�`�,5D#��`�u����2�)9��SͧW��*���sJ�!�0sɈ���#Պ�1<6�]�
�I�p��0-EJ>kF=�f�;}��EaZK�����׀f�ʞ�8�_���'�hY��c.Ð��8�w���6~XUg��}(�I��#����r����c�fvM�Ͱi,�S��l�PH��������ټ�,�X�3|��D$��8��7��T�-��yBb�/"C�?�W�+f��T	�����T�0˻�^�1]S����`�Uf���l��a�w��+M�>!�g�e_nG���B*��H�G���d�>��/muZ�/�K��/
�̒�b O�y�[��,W�rkX��uT�B���S�.t�ĭ�3^5ݟB��@��J� S ���UM��7W������6�;aT?~@l8U�odK|�����! M/]�����^��u�~V��M�Gp%���}�����|�(�GTsJ��٩-�nV#����Ա����	�*�E�]Fng��"Œ�p�⮌Z0�C�V�qAj�Z|8d��viRSf�+;�r�������a�8i%��i)�qf&��H t�P����TL�$j��m�ޜ��w��Hf|Q46�V�f!5(뼕��c'nl�V���$^�`�^'�]���ۖ�X?'�W�E���q�[���-EtV�q	����J�H��/b�,v�p����3��=�!����hi�VU�4Ŵ��A��۹\��ɲ�F�E �+��06�C��#�H�1���up��p��L��|FaM�}�+�S�����,5Z�������="��ň�"��~K1[��9j�c䠥���i�Q�a��<_�7ft�8,�|�5~��њ���g�h�F>YvI���ѡ�왅�&����#�	�1j����J�xn��������-�=��J����=A�P�;�p�u)e�5Z�[�`���@�Ծ?��H��/��Fg�}��.�MM����{��?d����&�D;AF���o���^j_���e�$��Bs�띩
SA* /�e9b�J�P�����ԚY��iT�]n����|ᥦ$�d���?.�4\��M�PsE�
��E�(Q6���aE,�������u����`yd�
���e��7
�c�`��>a@x9$*L��_��w"��i�sؓ�஫�@�]��+�p�|A��'���Ռ�8aHfX`���|�H�W��/��n.{&cX��]�X�`�N\k��vB(K�D��I�ģ�n�"�zeͭ�A͖E�k9�We��d\���7�%uh`�dp`�}����k���Ԅ�X��/�U��~0�m�z�E���'��Lϛi.�O��S��t�w��J[=;ks#pSi1�����Q[�^! $8��������+�/*��ʼ�Vu��H��U�F�gK��軠5���5,]����}T:���+��%_���;��-�n~_���WO����^���j�1&R�G��#�.W	 W�YdQ��)�[�c��&��B��|M��*RO ���1��#��y��l�j�e;Y����%v�@������w��!�	�hc���d9�+m�-�TW�x�zkR���E΢j�5(U�5�|i�DOy³q��6�QID�v�6꒿�h��!�M�T�,���l����*��sd��_��X�bJ�ٝ�)�vQ���`cf�M�}���Q�/�d8�+)�/]���hfi�zox�Ϥ�c,ą�]L�`A��&���|��5i+m�_��o���א�qZ�������J�����>w�I6��ؐ
1t�=O�l���������ۀ��Q��3IJ#�ӽ��\k�b����rRϲF����fλviȌp��gt���I�.E���!^���"�zt
�����g�w��@G��v#6q�V>������Iߍ{^��Δ�<����h��yŠM!������(Q��E}("�z�����L��q�lJ��'"�v0"G���gm�+�pC���;�jTx��G�N���}l�Y��w��2�0�;��RF�����;f6�S�G|����ٗ
��^�� ?y�̈<&����r��y���e2�U$���U_���4�*�
,xH ')_��N-� dՀ^��vg�����!]���=66K���]���A��n|�9т�R��	=p�8'Ѳޫt��W��jp��u�d*g�Qh�M��*d��42�n����쓌���
-��ܿ4�>
�"OIȆujp��/�+���@�eJ$?.����u�n��J?P����z�͚΋�ss�o���T���ٞ���k�����ބH|���4Þ�h�,�#��ynL�q��A�`E�A䛵ܪDUשZ�8#Y�z��O9��+d�N}3:�R�p�|y�O��G[۶�����<�B^>:��dxБ3�����HW���S�<|�^���<�-F]�SϨm������"Co9�����]���g�'!C����X�����o��=�AQ&^A���8�ޥ��}�pN{��Vo�� r��@I�c!���br��䬛K�6�H�cb@�NS>�?cոx}}�уh�]Z�vGk����^�)lk6w���!�5��2Ic�99w�u�@rU+�g)�< � ����fGu$dH��_#�Մ[��OP	��`�g$���?�Na�r�ƿ	of_d�bVu �M�:�lK�aKbMy��V��0U$ ��f]�¢ϡ��p�@���6!�V�>/1 
O!;u����?�vV�A�P��']pz+th	��5o��B��l�P�ސ��58{�=醻[1��(}���!l�@����cY�3k�	Q*�KK?��1�d�&`�g���F8���)��?���KP1� {��MR2���bIz���/�"+�ُY�����^�M�[Fo�{�AQ6�(�oi���e��B?��o>I���*)��.H��aΑ{(�=$BP�8**
����޹�ɖ!ݯ5��@�9�>}���}��,�X�y#��.qz�̧�OE���jI^��}?���x�Jb�Q���@�Q��Ĥy����Luj��?����NG����\��r�$1E���"�O"4:�>���'�q���k��C��z*�l�2S�����>*Sǐ�i��-]o/��$NE3ػ��7Ф�+5��2l�x�jy��EF��4�;܂D~�vf�W���呺K�ٚ!P	���H�A��U}į��G0�K*=��}k���$�x��V�y�KN���=�)�����X���%�5���;f�c�o����J����¿��z�N�����k�g9H�!��R�/��KqU]�3b��w&��Z����Р���X��d˿���s��Qo8.h�9�o�֩��"�!�}����k�v5��1d|ωEW�W����E�	q�!����l�ŀ�=�_��u�%�":��dh�������B%������Ym��>�/I�̀n�ݔ���4i	���+0����D�'*@�����%���gL,m��8��
����d�����t�f����į�cüe��	U;�إۀǲ~A���v
Kjդ��ɕF�G�F7f�ҏ�	a9D&��W��͑��@�O��+.5N#-����n᡼#�gQι��;iR&����9+���*#00y[~7�����<�)^��k�ޮ������d	W#�Ҭ���*�>�\�n h5}����i��m�|���Aؠ?�F�G��� ;���8ݲn���-˥����,U�,��w�����dj9���aai�P�N�&��2MC�������,E�����NxlA��HH�>�5[[)pz��)����w��m���g�4���&���%����eŞ��g&-t��6���������"�P���Ba|�D�'7N*0Ա���/��}���"�:r�Zo����^�a�
�@�E.]���ہ�ޏ g�}��^�M�O�����˹k���8fi�ܲ�O�5kY
�э�/�Y��F?<;(�դs�!�J����'�/q�:c-�>�:[?i�6i˯v�8t>�'��gs���Dn� �&��s��ڐY�k�|	����5�I��9�ɶ.;��,Ňo�S:�5-�뗹8].�goO��,�����^�<�ey��ړ����~�]���eYh�t��n���hj���/_��ez�9!��s7�A3�μ��{\���4��g�7R�xU��6k��\��V _���,�4SP���`�yȒ�b�\T:�K�W<�nI�IHD�3Y~r����ca힋�}(����TV������t
���~�P�P}�u���oa�W�O�ϰ t�<|�����5%?�5������%���}�M�k=�P�����m�+2��������i"�^�./V�'���؛���o��;�_��4�H������f����:�1�["�k1��X�{�s]_
�e�ۧ;AL'm.�$LN�I�[Am.QBK,i���mwҬՐ}��9�����M^��ꓜ�(t���}l�3 D�A���� �i�Ub��j�����}������ĝ��-c ����p�N�D�<����3<Zj:~���sϏ��?���E6Ndڎf��N��x)OK��4����7�k�o,�f�ŇG��"�ӿ��$w��	u��0.���}�Ԁ�q�����F��'�N��@Eb:+���](�������+�h�o
Y��Y��9���is�h�5|������k��NtR���ᡫ���^p�ʖ�*g���r` Ï��l��Td�ڈ� �` ڳWI����9
�(e������_�%��β�i_�����l���ƙn)#���`���
�|�#�!Ig�5���N�e��ޘ��qM�N�p�=$F���_j��2o_�M�/p���y�SFi�wԈ���u�q�c�ј�A�p;ӀR�S2pl�+L%@�:��.f�l#�����鮀�( ��iC�-��}��B5S������1%�ʲ�[�t1�`}|��q�WI��Y-3n�oI�hڿG�m��$R�kʪF������>?;�w�����sx*���%�(�u'��I%���S�R_�B*����{��4O�%ݘFmo-K��?�&���?���\-��-j���;�)��q)2E
RPh$:���:�Az���>���M4]��#�3(!֛�a���L�ՔH�V/�lu��y��bn�1�l��sS��\|��ac�{����\��c��1�RΆSU�uS�_��8蓎��r�)�A~�.�{��<�tn�}8�M*v>�T���P��<D%��s���](�:��̍�W�궰'D��ʢ���v{��SGT�#��Sm�EC�p�2 ���|.�B�w�(��Բ�)Sa�툩1R�/j�kQ��NF5Q h-#.N���� ��UE�U/��Kc�A7N�Ys'�
Ǖ����>�A�?�C�J��(DpL}��uʭ�t�;C�=6f1ss���$r\���wZW���(裒C|!���zm�I��v�F��y�dK5a�tiC�� ��Y�ﻹ�	;�rj�#�2[Jf�a�#$�ȧC&z�����o%hొsq0�{��/T��'.���~D������J�A<��a���?}��{�������<쉂�Ee�`y�*��-�e[9�b/M���߼۩n
}\��a%��OD�借V-{Euh�.UI��
� �6�R�<9w������H8c�,f����ɡg�3âUS-'�ZhpD��N��b~��!|��'�UZ��b��NQ�*�Cs���ΰ&B�*�ks, ��%oo6����a��M�ڣ��r��qc'�lgCRT��K�Ñ�v�"��?��S�d��X
 0?=����%J�#�g��a�y���'�!4򌋏w�uK�#^w����?fVFl+�,��H�J�^��.;G\ۂ�~�n�%y��@�y+>K2��{�ZX��m��`:�[1����樦�V��S)��w�����t]?�G^l����~�NS��S��sM�a$G���F��푢�pF}`M���t�[�Nٱ��k�Ț?b���BK"_a���ڡ�����|�s#i`�&.no
�~�4� j��"]_.zI�]`}��|���2���a~�h]�z�A���c��W��8�	ׯ$��T�F&���L�� ��V(�q�Q��Ӡ�`�?�&���f	��(^_d/lXe$�~���#q��>�h-Rd�ޠ�Q�R��<��5A����NYc�Gx)���V�O@���A�w1T�Ǟ*����.������߱�i_?�-3T��PD_�NU�������V������AfL��H�v���Xib�5 ���h,fۣo3"��bzFz^Ѡm�`9�	�"��Zؖ:{-�o��������G��&�BU�TƱ��ܷ͠}Õ�������d:��/�*�\neW���eL^�ĭmh�Jq��/�s{D�Hiz��v*<A��_W%v �A���ϐ�B3�j&D���;V�y��7�A���)�?P���/��|NtX��6u����
6l#���(�:��g��qX���ͯ�T�]�5�d��ύAQ�\� �Z4,sm��=��Ab7��R��j%�1�J���/�1���mAX��z��k?���t�F%_�'6�W��8�"��w���O9���ޞ�e�v{�����au^*͢���&��f�K���?1ahs�����렠ka[v������GJ��������2["S�/S����ݫJ�[L�����d��T]�ȭ�WU�0j���0�f�Z�'�H�lnņ\�����V^/1y�U�r�� [�%K'A��C,<�伥4�ew�c�U�k��A�7q��Z��䯷���T�c�V�y�
��.�;�h��#�P�J��I�4�z�܁�� ����qQ}���0�t#!ݠ�t���H#�Hw��4�]�4Jw�4 � �����}��f�ٱֳ�z����l�[{p���lek�!�_8����ym���Bq���,�"��vr�M�Q�|�U���Od�h\ҧ��Ӣ�̳7�*5�;dP����:�v׹�|od�|n�ž�e$�~�"�1�qw���H��>��j�#��J�s�E'��~T%}H/���56�/�=��2�����wL�_'}墄��C�F�ۨ�I�@���[�w��q��Nb���[��麱s���H�z���p��/{��&��P�09��Nx?[���J�6�� )�$O��#K=�M�C3P�r/�n��:�ov7��cc�n��CD��u��v�0�^>)��gm�&Ŧ�=��0�/��u���4�7���^����#����!�6U�،"k�DC5�8�8����I�s����^ƀ��-ػ�7V�zfxt�}#S����r�����=���ů�DSz�D.ũB]T���Z|Ư����Q����^R*��ׯ������������(��ӎ�3���\ˠ�r��MK����2�N��Z��>>�c����߆���l��~3 ��p%֩k�o*�s89���&��A
�̆6&E��f�s8���F�J<gvҫ20���;|u�Ə�����k[�$��8[�u��'��:܎���З�Tpq�o)��}'B��u4�8**}�#��b�����u)�����a�bG��u�t��Ѱ���B�7��mS~>�B�+��g���@:��j��f��=���ɋ�'���>_N|b|�Q�f6�V�R���9T������g�8u�f��u�t��o����'O�j�s,��q����jvJ��%���O�{?4M���W�k������n��f�Ƞ��}:�o*�?�b&s�)��0)�/����� �}�o���H,�o�Mi��Gj*(C����u#�|���qGQ��rb��E��:;��۟�'�juY���)��h�������'eN?�gw1L��-LE���E�ZVð�%����A�8K��1����b!%S3��+Q�ݔ ��:�ηmd�7��"l-���ty4���������Js�B��Sx��abj���djQ,��F�Ij���f�$Ks��P��~K��_�`�F��>wI4�����x��|���Xϛ�@�]}Ru%p�e0STTo��pC[�5���׫B+~������eyK�vrC��n��B���L7�m�z�E�[)�WAx~rQ8�b ӿ���}pHb�ѽ����(~���o�#?s�s�_����X4��8�x�A�3SS'(��(`{(��y$D��o�\������]Д�t�#k���+�Le!�}����V=������J52�J�p���"Ou�w�~�S�W�q&'K�(�܂����j
{u:q��+ݪ���?��f�=R�tN�b&%��<;�������쩮䣇�/i�|�٠Y�`,BV�S�\��4/����@�J�o�7&vr`�m_�[Tebϣ�#㊜�����B��Zm(���p�)c���P�L1"����o���4��{�c8��N舀���&��h�4��T��������
]ϳ�{?�H_-50����">��.��&�U�%���� V�.�A1������F��.8 �W�f+�� !�u��j��^�R���eښ1�CB��zDf�}�F�7����}�_#�h����(�?���,��u�W�)���?Û�i��ȁ�%��B����{X�
Y�kʝ����M	�*_�I�g"'C�WWX�
%H5���i�D��PɳP��dfs=[�v#�Q���V Gn�u$�ß�@�I@V߁� �B��t�C�V@�n��xN4�j�}�w��o�;�K� 쌖����L�uqr�^6}�sqX���u�C�8s⿴������Ž���d��N��}�V�v/0��]Q��!fX�8TB��y5	]��ytl]m���L$˳��_���v7}��A1\�MX��Np�SNNƹ]&�>Q�|�@i����L�cZ�qSTY4)�Q4��3|�5��ϛ���}�'����r�l��o��\���ڻ�ϡ�	젳WFS~�\a�Ls�#�q�ab.��DcVAe<�q��-��%I���,Y�z(��m΍<�wC��~v�˃ H���|�a�b��,�����|�D���"��=	g����_1�z�����ag�k�X�cI�q�w�����w���e2Ɵ��CP�.Pܗ���R:�:�] ػ��9g��lh�^���uݞ�����xξ�Yld*��5�$Y���%Q�p�����G����־� �%0Yy����P���_��#��d7��!e�["��<6/�����Q��A���~Z<��V�2,&��d���!�����}E���'���s̢EN���Ƥ���t �D\؈�n�8y���"d���>[�l��2TJ����T�c7����_��=�d���Ol����z\t�g�e�]�R�� F�E�{E����GZ�w�����*�%�qˌ��9�T}����9^������aR6᫠�Px�3|ZW�]¼�d��6���lзtx����[]��2�G��q���w�
���}�8��8M�	�:��Cs(Z�����J���������\�=͟�m��.�$(���|9�Y�8��yv"��$m��H�w�Tn��E~y�~�5w��~cGC�<.[k>�ٻhh��~D�h��'����T���K7�Wj3]~]��9���hr�W�D�kc�=|K#x:��S��N����,�Ԣ)����Z]��T�6�b�XҮz~�S��z�_�z0�P<�"ˍu���t��q�+T��HϾX�77+�ǿ����M�8��s��p���_]�=x����!j_��rr��/�fq�s�"MՋ8��:�A� 1���#��jƼBA.aj>���p�[;?�����B�y��
Yc|o�oWv��JH�	�����p@�*�����?�}p��?F�N��?U	 ģ
���13�w(�7�\�|�{I\}o��s�a��{?��9ϲTW�
:`{�d����b[�f�"�NN�{2���t�'5������;8�^�����iT�8�O����b����;����Yׯ;�9%�Xy�̫�GY�wa�����O�Tg�q������X�t����{�!X3�N����yyעZ^�Q���9H��R�ٍof64�
�&�T�ä�}N�q.���o�t��E�P��j˓a����n��6]:����yN|�f5�z���[u��[*�F�c��"����Otǳ�g�8��gOi݀W|���
�������:�<���&4����X��EV��!c��������R-�V��U����������e���1g.q����N�S;�uRW�nu����E�Tz�R�+�7Xܴ�����'���L�(xE�n��&���3�C/inGJ�A�����(��P�RGGez�~�60^ͭ��Q�[t.ѭ�b����Y�!�8B��r����	h:*���q݅�v��*�*Ǐ�)���j|��Fyu�9𯚼XDt<��ф�+���}�%��񚚍"��Η���;i����a"�i��O���ʹ�w���*��H�1~�ڬ�[Q���,�`l`s��"P<"ݲ�'�Uϲ�����FPβ�d��[���Λ1��Ie��^�O��o���]��/m�Rn� C� �����i��d�&���K��`,!��۝~ߕ���_x�7�D�s��Z�\�>�?��mj6]���贍|���ﺁ�̣�`����^p��{��q��s�IX�c�����!�ѿ#�˵�n��L���m�l�������j�ύ�K��� }���?w�f�(���� U�������F��IՇo;>z�/�jG
��eW�"�(�ē�+Ƿq�1�+,��-��{�v	��Ff��C����a��U�p��P���O3�2V	]���"��F�~Ss��?�x�?����䒛;�6��.L��ݡ1�f�*���*膾���oL}X�28PK�s���0?o�+�`�������d�K��XY������Cz!��8�������A<�nX���@=����*�kab�N=FW���3| Ō}�h�
]Y���>ɸ_?���S������b����V������Y��&x�˼���ۭ��u��ȏ �������Q��Ǭ�a�W��Bg7���s!�3��I�W�c�kc�8�+�Te<h�R�BcU��yd�Rfc}�c�$T�DK�4���l0i��g$�<]ot�G��*�.O}�x~�z5zo9D`�Ġ`�Y�5z���Vt��YԡÄn��Ir�M��1���t�����tZܮ�*���P
�������J�h����Uj���h�!��CL{�:^�C����gl���}��rSr9��N/N�i^HWc�RU�`�8T���龸��
PY���|T.d&7�a��.�΃oIÎ�3 �X4Pm�����>@�o7w�������$����,��.k?��`�Cl��AX�{�3�/l��ؤ��H��0���d-��xy��K����X<B/wް��7+ϧ!�sx/l�Y�L�����P���X'2���'���9�����JI��p�8��˻J��+D�pJ��A��Y=K2p�(��꠬�HX�I�#�[q��l�cܓ0@�?(D��E�П�����A��\Ā絥�����o���8�ź<߾O��c��}'���s�E��~V\�aɮ ��pd��7B���0E�P��O�;e!���'r@|�~����w�yQŏ�N��v4����I*h0>�4�
K?$�ȋ�Ր�eZ{�?$�;��9n2�(vDx�>����䭑f�s��t�`�Q�:Fq(������������d(���������	�cH��W����3)�X8_�7T�ܧ�,AIP� �:���j?a��� ���
`����S��I��"���)(����xe4��|����D$L�n��wn�Y%�����-|�i��\Ďވ�&�P<��`�[d~]{'�گ��1Y�"HY4xm��N�/h%ǁ�o/��.Y�㓲��,��L��Y���3G����Z�Z�2~0Alv��u�9�vlņ����`G8�G���zI6C�b�����{�K�?��Q�[qb��mz+�Ĭ)��?��aq/<�ä���X���I� �{g�h��z��Y�wD���V�w�g@��P})+�l�|a�l����� S��@p����uL�� �������"�뺁 �6��7�jN�K^c뀂W�f�Y��%Zl�2��R��jk��r����<��.I���*�-�Z�@y�d���I(�n{L�|d�8g%�[L����C܁�Ip�/T%Z���NM��2N8�K,�h<�W%��|u���I����â�E��;�/�,.�&�
L���S����t��.���@99q���̡��9�nIgN�Ӷ\�K�'h���kT:)�����#z���������?�g(����et���e[��O+�q����|�.d$�52A7�C�5�z�/�n10�����`���v[2�u�Gm�?W�uu\��E��"�+5��ÜBI�rK��~4���H*�)���J�W)E_نT��
�$�D��$�KF1���������m�))�xq 0~����ĭ���oC���z�* �>��(#i��i��,�~��.���p+��N��#���b2]�OL?�����ʍ�2����G�G_�o��]����mkB������m�%�4"�T[����u}-���YuR������9��
)഍}��[N�2�Mƀ�ˡ��~K�7lN|������7)Rh���Z��d�Ϟ�69cX��'+�)::8���'��y�We��*�������핀�j�Yν@�jYt5����Ǐ{*hG�f��EN:�Sn��ޗOQ}����;��;>1�#O[Ky�hR�G	�]�}T��d��v*�7G�y��z�BC�s�3!f�-�{)�xҏ�tL�@-��Q���bO�}n���.���~u��8������eaw�٧o�Y˾z�2\((����u���Q:*�4�4�y�ʴ�k@�ǲ��`:��q��R,�����I�n��ص������^�1��έ^�bd�
�I�2�~ms��Q�JYN!�Pe�ʋ��A?/>�;tT��S(?���t	5�����9	A�i⎫�(��Z��W�㠒�ā�Y&f��A�`�Ш�LM��P>/�j���qU�m�� �7E=ڭ�>�6C���i��2��=j՜�+�"d��vb�-�B�
i7�=���1�l@s�o>T�y*"e��Sr��!�wjf$%����O��Zu�#ֿu.G�Z�WYC|�|��%��C�����U
&�w���*��&Сe��tn��}�E��	��R:�-ɗ	*�yK���������'� �/Ǜr����L���#R
O�����e�˝��g�r����ٓ�T�W��'˕2����F�B3y#�ux&�M5(6q2��r����*���F�˂̡dn�d��3ˬ�6�� �����I�W�N�����0���M�h���5qr�M�:J�'���瓙�P�)�4{���=l�t1���&���Ԩ�H/�����/�]�,�������a5Gp�@�����j��zꢲf���G���� H�|H���ӛ�	�~2��5�ɺb�wn)��(��
#�륈�S.�6�>^��n���(u������kt+}��M���,>
����,(�{9��7�K�YW>����ײ�Z���):�)�W��q�5�L{�`Gw|F�X�E�<��yY���=�L"1����aR�m����a2J'�����Su�f�/a�=�c�-�q���{�� +7�_��.B5�7W��@]���G��ǡ@�O �ON�Ĥ����'����I�����9�V����C�Q�-�-� �������0�v
�Sֻ�q�����˪����J	��c�f�!�J�-N��`����v��I������&�1�'���
�M���{�{��]�o{Ȑ2� 
��N��E�Y��t$��x�N��<�A����M���/�ػ�L��>�ɑ!J�n:�--e�rm�3�O����C��y=H ���jdR�ϻM�9_���KMf�k��i���I3�V�p���r��p��D�ߡX�\Q4���kOYY�r࿝�bZ��F�lU�i�8����9;��.BU��[�$ w�42W�٪�&�+�s�J��#�X�������f�/��* �UC����Z,U�5>�1�w�n0^�O����[:*=M�5\h"m��J�e��++%��t���t1џ��d�\S�ȅ�
4�ԛ�`5Nb�G��LP5bw�������{	Ǜ Y�+���q��W>�ш�Ox��t���\�d&�.�ۦF�iab�dy.$��B&m#�*��q�b���3�2 Ќ��G7��AObȝ#(-X�3��hGt�UU=�n�r�ƀ�����_ޠ�ℨV>���v�ة�[J��)� �-�_˰7�q���F���L�2�r8��jd����3S#���	6�J)тC���?~����2���ڱ���W�ŕ�ߟ- �M�vQ�-�$�k"���dc���V�ˍP�q\7���a4g���ptk�8_KX��6_[�8e(1�/,ԙs�p�BB'�_��g��ǡ� ��c-��f	E�A�� �@q�t�&��6*f���vq�鏌�����lن���У3����{�A���
,�aG7�:�2�/|������Z��ZR9��C͋�����êO8�X�K<A���Fp������,�����5P��V+'���(O&�bNhP�d�6�@�o� �y6o�-��iD��"��{�-E��\r ���ع�FHe���O>|�טG2���s�D>_�u\�_��A�,^��n��ĵ!ff=���b����;ۮ� ��ۯ���P��Cž�WӮ�Jt�	�R[��e2�]�_����h�WU��6+B6}�<S):�m���J�2�?�>��A�ؙMp巣��D�)f��������&I�ר5}�h}Xnu����G��ߣ@.�(7x	�4���'��p�:t�_��q݀�4D�`ڕ�(����RW;d�̌�yX���hX�ZUP4����S��)ftY�4W�Q:��ר��z��"O٢��foo�����y̤c��
CW. �����!_
�+��j&����MΠo!ؖ%��Í;xE;�&3�>�Q�e�II���>Wi�Y\Q?��μcukS��es�wS���z-6��A�g/9�d��N8zd�~hٽ�xx��@���@�(�/��P* ���\���QWWd�(D���jХo���ػ��ms;�����A�����/�98t/�b3��Sy��E��jo� 05�AJ��l~���okuH������p*o�سﲜCc�1˹����ǿ#W3Ks	�"׳0ww�j9���&r�B���hݚ�D����Ԓ��C��"i{m���ˈsYlW��d�N4_�9��KqX,�x�49"B5����N_ʹE}�c�b� ~�#K��C�RU��w��
W!�x��p%=�9B<�a~��r�v0Z��29ۀ��ER����F����
�؃��4,���ߺ����kKx �ŧ�$H-@0ݎ��܈����=�����nFO�A���d���7\?j��y�
��8�̆��`�H��������M�@���m 0jd�@��	���� �����ueE|���ĝ@��!*C�H���'C���q�a󱽃l�V ��he�j�E��Y�*Gc)�.#�?X�O ����"J�R#�߶(�K���FT�/҉pOS�t#)K�T�����l�I'�WY7D��x�iC��M���>]!���P���z�1g��4y��!u2::࿍��<ko���`��l4��
I��d1�0Y�c�S��(�\�J���W@�@
3� ��'��^�k�PßX���X( 74����f��N'�ۍ5����L����:\LN�j��X�rYQ1>�^MJ��~�F/�֏P�L��kj��C2C��EA��m^5��q~���!����a����Z���ӕ��斥<SD-�f?�r�nZ�7��94]�B\:�2R��,k >3�!$T���@KX��3,���R��p�����0�m�:��fK��c�Y�����B��0�^��x#�!�!V�_��M7�|eQ}n�w;|5���kr�\�|�x��JAE�C�k	�C�:9d��Ԟ����I��x0�B �,���vÆ�sX?�Y�Y�v���O�f]����:=/l�x��:������;��V8E�S]�j6�W���y�̈�F,O���+�J���B��F����C������p�E�B]��$⢎K-�Bw�*j���I�YUJxK�����K�x�5����;���|�ߤ�M���ݜm?I��l��KԝCp�X��l���L�*@�����e�楎*�l���QPsl���_��;G2�'6C!�w�|i��շ�x؃��%6o~��MS|��m;�J(�D�H�!���B�m���W+�\�Tf��Amw��K�2��|�������"e�,VB���i=T�G�%�J	4b$���2���@�u�)�_�4��9t$�x��K�C�ZJ��+b��?w�pb����wI<-�*�	Ke�#;�U�]֡��	(0?2�a�i;W<j:�X���b�+�t���e(���i�GC`>�m�$z��<V�su���ܬ|�w�L �/|�>�6�&h�8:Ė��qP΃������1*���(�0cx��K$%���%s�N,��xHR0K���z��X@c%��O��LB:�%���(����f�>����Dbe-S��(y�?TN��!?� H��_��r�}$�Lg��B7��A�-�F�uW
���Ǩq�@;
̶�� G��j���W�&4s)r!�SiL��	a�M�U�k6C!�9�9�O�/#�ҫ1�Rś�{b_t����y�ʡ����C {�;?YTZ��Kc��!�	�/&�5�x��+���6�k' ��{���*B�Cr�ρw ����:C@4O����iI���yȎ�Js�"�c#�Ɏ��
��r˻����2�����M��_}�j�cP,�/�M�J�IH+�G\�\՗С�YF�R8_V@t���uE�O��eD<6��'x]+�d��,�&Yp�x+P�fN�̡��}�{�{����&$��,>�����ǋ(.C=J��|y�c�y�?�(��eu� W���4͑��	�<	9�����1i.����������_7t����uYZ�׋thG�}�&ȝ� i�RO�y,ܜ�����~��E��y�F�/,���K\�.�������Lڀ��A?VJ�W,P��ሴ���� Pk�T��uH�(&`���2h�cCH����w���(��N$�	F�������H"�n����2k�|=��u��j	�����fT^r����w_����%`�������P�WL�@m9f1��ͪ�G���m�u+��EE7�,�T0O�]�Z�v�`���i�~�|C )0b��!��0|�" �o�ʡN�R�,��aM�p:\�O�������p��\���$��q���1:�m3=_C��Vg�����  /9�'z=� �	�=_@
�0 $�]_�,*�6��eQX�K�^I��������dYol�:]�9��������8D��,~�G���3��S�ϊZ��q@|�0Q� ���}t���Q�����/m���r�uv%B�ri�>nB��� D�ģ�6ߢ�@N�o�s�f��MK]ث�#?��7*ʱ��y<���I�0��0��·�;�㆐�|� �����,��^@UC3U��4gn��K`�*��Y( ������y��x#1HtAUbAԔ�&�q�{m�8(<�{sH���5����a�ׯG	�D�e IUy�<�NP�q_�^���zZ
j��/�UV�[�٘L^,�윓)���3S�8>�Q���T|�0tEw�V>*nj
���iL�N}�2�ɿI�gL�����E4��	ȩ%,~�3(Z�bR��/��B;���X����\
c�͍�#��H/��?&��B���;�4.ĺא�`�,�s�!h���@���W�o����׾�c��Bѧ��F��C��Ƌ���ۼ�$K+uAo�}��įtA�#6;<!?������	���o�!���$�t�B�)w�'6��z��ɏ��R2`�UM�b,A0%�@������nҋ��>��Ht�r�NwԀh06q�:�r"�Y���)P��Yqk�\1����>��=�X����.D�����\v _��кɑݻ�]��
+�#.�pǛ�51S�u�S娴P"9%1��m����P'��&i� vv�Y�`C�R$ 'W.l,C���w,��hu�g�>��4RgpS��bu=�"�
�8[X��c�x+��ڸ��*Ǥ%fl�vK�* ��r_߉E�c�2����=��h���
��kni�'Y�'6�|/�&\x�����+��];i��}�|M䷧�aȑ�t�n\�=3��CX�.��� up��(<��:�@g���IigjP�ͳ�������ʟ`, ��	ts���8&��w.����K�a	ͬ����g��YGG�O$�p68����r��k���C�*=59��;��sL�c_c��e	��x8?/�����:[@��^�a�$ht��HS�cN�o�����#6�&�h'�\���?F�c#7a���}���n �{C��+���^�(�r�X ���h콻!��!���B6v󓞟��<svAy.���-Klդ���!��β�����O���p�{6{D>͗Υm��3�|���YAq��Ȣ�P�uD��i�Ħ^B�A��\��- �)�|�'Zl���uL����@���p�t8B�/n#�b��x�(M��r�YOd[��KS#��1���۳�i��ށ�-r,$%hw��Ԥ7!����F��Ua��G��~��S����!kEK-��!��B�-! ͆�X��RM�گT��l�; �h�`��ի��k�n��K�榧q�v*�ʰ��)S��W�W¥,�����ީ�|aw� q�sٰ��t� R<�e�V���yy�s��|P���5{
H?�����%V*�1-�U�JJi[��*M到�x��c�Θ�ʕ������|�x�'�S��o	�7���YM��s����kf��j� �H�]l�3��C��+�1�����j����������G-��}	L]��!���J�2��/"�6�KE|1W��ũ�G��"�-����%�3$V�G�.���-y��D	�y���CѦ7���xd4k �ۈ7t��w��
��+�G��(G-fi�/�f���@���H��G
� R2��h5��9 ��6P7P��Ѐo����m'~���W$$)�u��
�D�0vU�ý�9�yj�g�r�wO� )Eac�?�>�Xߑ��shf���
�K��J�u� �pM~f���j�'ɫB=rX�4�s"��u�|K�e�����k�S}�F$�+�����aE'f%e��y�'�S����4^<�\����t�|=��p�G�=q�"=���S�?զr"�E�IC�dq����9@�M�mUkO�ԹM뺕�B{���H�:�L��n�Ef���e�����_�5)	�F�d�?��C�gD,]��Ƕ6�tVw���[���6��������H�$�oX�r�qI`���ç.e�Ʋ挍-�w_9���;�^M�Lifa�/�i�#nRH�-����ѓ��A�[���J�^kC$�]�
=�7YWLUӘ�a��oe�b�\KE�h�l
��jV7��(gV~"n��Rn��W�H�ֶE
چ_2+)���Ij/��K���t���Y�\����Sg=���|�.���+�է.ٚZ�7k�0A/� -4�i�mV2,":_�������Ɗ��kf|�*qw1�y�:�r,��v��ݔ\��}�P����g)Hj�8y�6^�e�-f�9:��P�vR:����@����hQ �_ډ���4�Ц���Aj&ס?E�e�j"U�;џ����e^�`2��8�*b�Z˱�$V
���K[�C���!��>�ޤ �+7ܿ�Y!=�P1�:��{c`���ݭ�]}��[B5��H�v��ԇ�t_�D��@�lQJn��ŭ
��R�Z�����W�H���-���OVU�֡����BPU`d�|z����8(���0p!/��ͫ%��a�T��af�Ӹ���aW�����x
���ul	��l��&��z�7ӏ��*����k��%!Dk��|��b�v<o5��M���e%���}��|�&Q���>6��ئ���@zM���\�x�ݞ�9��(��,�ߦ��]e� wц^�D?o��c�v�Ґ��h�k"P/�7�v����������X��)�D��7��tm����U�˩�|Ǒg£�%V��T�}LT�xB Am��G�-�s�
t�:a!�$��N�Q5����c�$�c�a��'�3vx�_���͹e_�B&a���>�<߶ P;52+iL�ׅ�N�:�;�J�������%;��������ZNn�c=���3���i(�� ����� �E�{ns�K׿�Y(g=��3�|�X��;tK�ǡǪ��<ou1��ܟO"���][������l���G*X|��pZl����]���z��Xq�N�ٗ��%U�?ۨ��W(��ܨK�k�`~3��6�czI�f�?5�^�튮:�4�v��9`�h������{����C�d�g��+-�yB�\�N�`D-.�>�Q���D����TKKc�� d��H�Q��n��3�Tc��R�r��}���u��h��ݗ$�P���V���?�ڝ��w��ɭ�Y\��h����V}���������P��"�
<;pq�4�<�#s�G�~�U;xMqҁ����]޵X'��{�*�����5�f<&��ӳ�.�{D�ߕ-?��@�9���n�$<�<�4!(I$؄��XSS���<�	R��R��B����rX{×���9H��츊	�������{/��Gh�@M�T�cN�X|�@aߴ�����	��Z�{��L�?�0�O9�+{ɟ�Oph�)p	���h_�bj���2ϜȠyab���c�)S�L����+�SK��V�Ч����;������)��%�z���#��5_D�l{TWk�g�G�罉������e�.u�i)qKQ=h��3�.F�@c�Y�[t�O~J�R=���4\�=�~z�J�x���� �Ϊ!����֔�e+3o�˃�`��͍Q:��\�9�^��2 ҂j�vZ,h�(S�� :La**�>0�8�#�D�nn7SD���Ֆhq? ��,�&��,�����?A�W��,��K�i���km��n(�)�L��ğo�68�KP?��+�Lݨ#t�*�yv�d�3��d�oʫ��5�]���V|���(gbJ�!b����?�d�$��b�.�^�$�;��Moj���C���퓝 �pLr�r��%�3�6�L��� \��,�n5��h����]���>6�d#��%�>�3��+��W�;��O|j�R}�4��[.8�bO(rӺj����S[N��t��O�M*rs�ʖ'"��Y��[���%WSD(��uocqg�L��THP��ia$3���ֱ݃BI�n��H!^�㮓$HI����iP�$��sBx��{1����{ϛ������}��gR���k���7����ti����N�X�� v����3��@��������E$��e����Ԇ#zY��=
�8܏d���[
�?�D��mY&��dD��4��ob�ί����rHx��aC~ӯ|Sw�eq1�~Yg>��uMy��׾�,��lI/�6f�G���I�Gdw�����z^����w��mM�r��T74���u>�}�o��	���X����Z�9�SǪq���V  � �cj���;dqݕ�g����q�hA�K�`�\����i �Q�V�;�������04d�X]/��I9�x�ZK�w�	����&��@�k��$�>8���P���;�{��b���8����0��+B�.�`�<_�I��}�{�9O���7Y³�/�8A��u��)�p����2[�|ۛ�A�Vɒ)z�SL�<�;�� N�G(1rp`��8����Z_�jw��*Y4i'���Y3j:��/��$�-�#*�� ��M#��޿0��7��[����)��W)O�h2�|n~0�|��Q������R�^r1�~79�,g��O	�ykVL'��c�ύ%#A�	z0vF�Iix�392�κ��W�;M�d9���4fHX�x����Ɲ���L��9�q���F���v$CSO�+�����;3K�6X^O�v�ӷ���E�b��א��8�աc�OOlVϭI�,�	'C�5��߇J��2(���e�͞��:_�r��l؇�I�Qg��,�3 ]J=���
��UƏ<��xټ�f�IJ����R�d7��9ږ���h{��δ$�SdK��<�*�"�S"�A\�e򛂖/�3^ h��+:�6��#u�㾱�y��m#��V��Ұs��?mlsv �t>sQ�՚F�ޗX�/7�;�P�<>�w�	��e�&��H%{/������(��B�__X:��ಌ��0��xȕ$�cI����bJ�z����Ç3�k ?}�[�@΢P���fe�?�*�@���R�Gw�.e��RE@�(��f��9�S̻W1���}y�Y
Q�xp�:���:ڌ�_�m�'��_^�i����Ѫ!��n�[6��?�
��H�j4��5�?�� |����7,}�ʡ�ћ���E�or?<2�����SQ�=$	���.�cT{�{�~�X@Z��Q�)���E�-dO���X%��x�W��<���n0p�$7�c(?��c�����}`�M�_^���Y{ �ɲ�V����֔��V�c�[����%�]cM���7��U\^&rZ�><��X�$��V6~�k�m�{���I:L@f������V���	JC[[x��B9��7-�q)+����g��;�PƊ� l{3��^�yo���m�!��8�Ɵ|v<�4 ĭ(���*Wߑ�dnT��Lf���5��++.�����oR��:�þʢn���0l��[���͏�/V���w���6gx�m�	&��y�[����k���>�g��a�������D�1Ϊ�0�?�j��n�Qf�w3�ʮ��!2%Xէ$��2 N�$X,�����[G܍�W粆��#��o��J�ܶ��Fv�R6UE%�3��<����0e����m�y�U�Y���P���@�{�!{�z:N�@F�9g�H=����;�]���(<�����N�Ge4bQ�I�����5�/�H�ۘ��A��Q�h��@+�T��v��wE��f�5��-S(�`��r0����8�$J�%��!�*���S\M�5:�{pww�w��\�݂$�;�݃Kp�!��������?�V�S�JR3�{�����9ӃG=|� ��q� :�NǛ����Fc0�f��>$9#J_䪼� ����9�jғo�M[H[�L���>ETs��Q�~> l,-���/d` ����"�oкՂ�,4���#�>9~� �Ȩ��mк�6�ҶF{[��K[�/��G���ɭ��&+�N�E��yL#F��r���R݉'4��&�j���}iz���sił���3�G�. vѯ�?!�����Bf���Z��{W�����z���:Y�t���p7A����z�1�8�&ǩ��t{c
�U��g
���.16�0��Ve�����4wH ��#O~��u���F�k��ل?����p�g���1�՜�_$!_�?`���6���[-x��d�z�ST(��%^U�9�&�Lw��Q��1�����&�:*=����������WO��exPv�l��ޗ�CT���xs�op7򴞝�U����M�x�~�z1�����JXFދb�'����Z$�t�=�`]�}RwG/�;��>o-���)ԠyY{�]�LY���ވ�R=\�0ZKV�{mkί�o'�c$6"|YJG�V��[��Nb�L��B�sV�����˿5[7�E_�G�`B؟io�(���~n�;Ǥ� Y�'���~�Wѩ��֒u�R�|��i띔�D(h��C3��/O"D�A��ƀ�5�Q�PzS)�`��	�<��\!�K�p���^�m� �Sv��ń�^g�N:#F
�jy��;W�%�q���X8�&#G�@x�F֖ݟ�O�Xx�V~Ub$�h�z-I"�$?{}�x4qLˎY�IC���̪A�h��<���ѝ���	��q������i��2`B�h�1&ˎ�笖?u�*�E��!*�Bd���J�W%��ʬ���=����lR_��ڴd)��~{��!��u} ����S�ma7Tj�́<�F��d��l���IOJ̄����;�6�:��Q��,��S��Uo��<�6�~�	L�{J������UI�g˷�qId��_п�¼'��`)�����!�u�K5V<i�����m�!n�������J�ۛ:�(�.=_�G*8��E����rj<Z�5���6xr��iNѠt�SҪ�����&��~֪���{�F�P���Ni�Ռ�^�G���Y�ӪD��r�z!� ����D$8I��Q��mKY�N�-�B��ā�V��\$�<9�̫_��C-T�5�'�BYao�޻�͸}^��x�{Pw}�*}�t�T���N�L���Z�����E���*m�7�����ᤵN�)w&����{�}��;fU����6�%\��9\6�Dt���b����j-�.:�2�V��P�F������<g����)�A�!\����ϔN�\���`ժ뢥���4:�9��G����/JbD�cbH�&P��W���D	Ŗ���JJ�\�F�F�I��-Z����J��I�k f;�Mo��>!y�`���TLf�>'�94h�lP������E;��gT�"yf���J�z�/����)�N�du�7�����;�YFX~��R�҈���4&��nq��T!3smv&zf�����:ܾ>�lJ��JEc���<s\���<'�����H���xc�
s
�Tm��$X�0D��;���&�Vs��?��$%�lV:a&����>sb=��=z�D#�Yj:�d+�S�o�~���3��;�,C�"b
�]|x��e蒗���%�� EƂY���	>Y���a�e�Ņd�6����7�g�^#_�����t��m��[M�Q=���A��	zOe���4�V_T���3{�i��4wC��Z�"э@`_
�Y0�tur��?Y�<Y�֖g�L����zy9I$��/��F�9�����d����%lxNo�=����W�T�M�ǎ���h�1��@ҨR_��f	�61����y���=-�?�&��rV�h��*�K�:�,�^?|M2�mM�� �V9v��ѫ�*`Dr�������yz��Y.�Y�W��x�&��9�w�0K�ռ2\w�nH4q�Y��
$'����(Z�V�"QG��2Z�5Ԕ��O4Hw�x^��LZ��I\JRz$VR��:�����&���������]�����qfT�(��$H�Uڤ!rн7�A�X�Q�۷+�����Rj�đ��>��H~Z��e�`��<`X 9%�~��? ɾg*���S��H�*w]J�ND���I����'�m�)��A9ip��JL�h�Ĉ�����%>�y@@:�4/���r3@	���\+D�-�D[y��溉;���Ut�9Żp0ɵ��R�A�S��ʠY�����]k�ߍ���w��.�,Wä��g�ǚ{~=����Tۃ���h՜�>L1��.��B�l`$��5D~L��F �w��)]z�3/Q�����\��*
$2�n�*q5(�4S���|�2�Q���SX<���
@g�OU_������9�����G1o�wp�u�&iC}�ar�b���L�wT�1�Ñ���t��ް��c%O�~)���x�>����s�F%�*�uĹ�	��(���=��}I�MFy��Jͬ�A*�,W?�����-]��$��'�$�l���k �e]J�1�rVl��w ���a&f���ǃQ��d+Wĉ[�V�ɽ��:j_�������}���x�"���ϒa��F�48�Л�"Lv�6ō(!��������}-<��,�×������3&l
�j����OY��0��o枾�iYSY���hm����uѦ��G|�1�+�1�A��y���Gg.���,��N��=c�S4PP�1�3I�����ͥ蒡�]�r;� ��z̲�4�uF{�~Z*܀b�np�"P<'���'��R����e��	P��O8������W˃N뜺����ä���Q���_��m�7�#�lf|�&v	I�%����Z����)��N�!��sn�D�rS����Z,��"��:?�`j bh�k}RL��>��b�&������mj��sy���9�z,�"+�7���12,�K��-@�ϤM��Ҭ�
�bx�%�W� ��P.��4��=�؏��@I���Ь�x(-��眄[6��F2+����Q8����YaAlC�\�L\"�=/�w9���Ttdz�ɉN� ���Ҥ��4.{1J���'w=_���5E���Nw<!��f����G�k�j!���2ǒ
�Ӹ4Z�_(�]N��
 G��+QN���y�X�O�!�\�2V#5N&_�іo�0 |�NEl��Y��4�$��!�*��
�b	3�����P��G�v��_�!��͵tA���/�/�y���k^��:
%�T�J��.�h�z��Xڄ�#\�U�7�i�ʵ����J ��m@���U�e	���n�I��;���z�}*��s$�º�La)��� ���|ǩ�#@z:x��}�ϸcZ��LB�Z��iZ��2D̉�^L
hOd���b$�
����HU#����d�tW�.�4���ezسY���I:����S���ضke�(��a/���1oj�]XV��g-K�_ِ|���D*�Ts� G��f���Ӭ����_��'�֫#O�za���.�h�|)�0Qr�g�K��Yx�E�ӖVd;Y�s`�aRhA����AZ�c;ЮV�#eD�o�J�+�|zʨ��Ө����*�3*N����L��=���Բf�aY��نɋ����Z趣,�ɥ��OMȁZd��m���c����tBׯ�F��p����Y�q���z�(wV�O^���+���Xޣ0˖=��z��g���6>J֮`9��E�qU  M�E
?�I�2��yO�T���m���(� ��r`gk)�Y�H�j���ȳlB��^`q�y_��ih�-WCa�A�	�z�qav�*���qj��v�DS��Ng�h$�� F_��^��6���r1tvtY�	P�3�	�z8�{�
�ś�c�q���ì�(�\�=T\A��t��O�L��?�d���?R[�3@Ub��)��R<�S0�(����%�g���Y���IC*i�lד�Z�V�Q����5I͌U>}��9/4�#�l�c]jl�{��%34�P^�E��u�����cY�V���a%�ƃ?��8��'�RF�;Яi�^/º�m�zg]�Ty.h�sb#�J�Ԝ�w��d5�>��uka�O�I\�崂���ia�4]kζ�'t�%��A�r=���(mX�	�ș�o�0��7&��(սb[�� 8���0Å�o���|2��8w��=��)kD��I�ŋ�d�����I#+��ݽ��e�����k	�͏�@ar6U�a��x�ìv����iC�� _.;�9(n��Y�ʧp]��Οk�����6kPh�"���V���:/Z��i�km�G!P3XX�C+�{�Ї`ghh~�d9�
a��%�q���?NR%W���1;8���%��A�����W��������x�e�@�C(��k�a�+��+����d|F�f�LO����Pg7}���-��èF/�FF�_Ү����nis�9QY�f��M|��� ���Za��G{����4����y&C�kmM��4�gF�iZ̮�k�V�Ƌ��7��X�4�������	J#¿C�������1����:�Y�<��P�7��O9���׺I�9(C�0���vF��
��$�}�8y.�����3?3��٠,�ph�Y=-IrԳ�5Z2\�#���6����>�����{��#Ɏ_ln�@�R����h3�?���_��[l}�X$9�������o��=מJ(˔7^2�>m��/��ԿV"I|gv~/@z�? ��ME�b���h�"t��P<���`y����ꃊ�w���e��R.���ŷdmkd��  �&���.�	'
2�b���L�{ꌧ�Y���L�7�(�ZpX��%����p�������f!����a�����O�/�����8�h�ߘ�Ja�|�ʗʷ��s�t�f�܅j^X�)y������NHr�<h2�!�w�+b(LDG�%�{Y͔[��~�p�\�2_�:%�E��r�S��lQ7*zC�B�����&�^��G����q����0�Fz��7�F)w��0l�GY`���z�R�@_�M�0�S;�����5Kȣ:�òtK��;�h<0�Y�S,�U ��(�x��P�&W����>r�mVE�ᨖe��f�;_���Y�.1�����R1A���l���G���|�as���[���h|�(�ը��܇�\׎��s�sB�9�]�\bS�l0pWf{�}��"� dF{�G�]\���~�N��#c�����Q���e��*��z��w���D5uE��f]=�W���6�9Y{�jo@C�8����������)з�:jg΀U�;��٫�î�
���ӈ=F����$.� �Eq��[�������ˬ=��0<��O�&��-�׳��7��w�z<XI�������:�@�Cݠ\KO����:���b�g����QO��c�8=@1�Š�.�H�[["ӧ\�����Xq]\&��w��Zw��7U&�����^0�xK0�'<�c�g��0*T��,�9��ݛ�P�4Σ��"玺���(�"�'�f/0Ѽ��M�B��p4��<���iR�����
�a���ﰝ$%�Q��.4���*�3�H��/?�ԄI���5�y
<��!�֕�;F�4���D�,A��FK'B'��S-�������>�ǁ��韗�T+����t)=V�S(G]	ͮ��+���4p��֐nB�X������n}ģ�5�J�Y���$E�������}�4����D�t�Mo̪5.��o�	l+/m4�)�����*�o����Y��P�'��$dJ�M��	�e�jN�x9ܝ=�|�QB��zQa�˂LL������c1��O�����`H�-|Ș:���p5�������}(���V��<o���D��@�n�|l�ykRв�bz��[
��'ʹi�=I^I��HV��J�ne�9y'r4�ލT�D�D�h���a<p�[Zz��Me��Q����]��{�O:��NφEX��ʺ��Yǂ����Ig���N�T�'��?V��������=��0A�;I��!U�{���/�^�d���2��r��	[���<���G�U@�i�A_;s�EyrVh��k^K��x`�?����:JF�:P~m8��`0��u��d�/8�a�ۨS�&@㫞���F����7��r��d�^�bҴ�!�,�3V�	!�w�
U�B!SL9��p��`��a�����i|��]���v�ߛ�P7�%�B���d�ϐ���s�A�8�c=�Y��ň�]:ģ3/�&o��0,�|�5�_�x��1h���<��+j�؅͠�,o�-��B���cC2N�B,���%�)ȅ��p�����FOv�s�:G.���I\�phYH�f2v�0��D�W�l�V��Mq�`؏ߍ$�n�/�W��>i���	�ϫ���R�?z��؜�[/�gx��ġ�v*�:ѐ�Y�k!t��B����u���l˖�h�s�5b�F�J��*ҟ�i��g|��c��ײ��Z��h~�<�<�;�����1�[�m4T83�""�h�i�'�#�{GW;�����G:�+mZ V��T�����׻]3	��ĺTZ�N�2�d"F&T�S���1��� ���r���=c��xQ��d|��i�z��hGt��Hd���V�M���l�հ���������K��C�.c�C�T��0��Yy�6R.��$����&��Bs�D�Z_��"��ڐ��)3;廉o,PS���T =�	 'L�.�k�Ǧ��:��\t�v�V�Hg/G.��ځ�&/�h��� ����J����`xQ9�F++<�xc�{��懎{�ጓ�!���=��u�ߋ�����,�Gl���CM���L�m�5G���q�m����`�Ţ6�He1A�I�6U��@p �j��/��MV���G�c����N�1�h����)%��9�no�coR]���@�xR���\��j��}޳��rW#e8����z�W=o�6�Y'�����[`N��P�x~xI�����Y]-G:O�~u�_Lm�o�Xќ�b��������	���
����P2���������\3�<#S�Jj��d�EyC{ĊwW��'K���e������(��?���V ��/]]u��v��ygy]�'���O*����q;#Qv���'���]����d�v(���g f�>��"�[�ל��!��d�l1��d[e�&�OQ�
�g[Ggm��T�(����̹~��;��cf�GO���-8��a���w��(6����_,����R�<�P�a�<��d��Qn�=�@&3�G5+}�2�B�n��Fط� @凮\\��U��!1b	8CUd��Oa�|.<<8A��o���q�(��\�:\^��>$���|]��N��qSqq��#s}�PP�x.+�b|�~3G����KA��+Z�G/w6��B�CR���&��d�}O$�Ǧ�i(�z�@��F�V�b)�'�i�C��*�������F�j"�:�!(!f@a\�1��O�) t54R�B��B��,{nB�u���3�/�t�2�gǐچ����z�@�:��=<|�k��{�SL*C��uz�l<��d��ly���y.�Oٽ�&�GL�gm��@f��p�Z�b��&a�؉K!��JʕB�\!8|MTG��-w��w�(�`rm҂�_wk���A1hb_�WP�����'��3��O�GMt����>�@����;��*f~d�g�j���P�-�Xҩ}s�M-&��@����$̠��4L�Z>����G���[������H#2f���f/܃�r)��THuH����H��<�:pzT��[���XVRd�NIm�6�Y<E5+����s�U��f���Ay';���l��H)
&����\p%��L6o��F֩����m~sd�Ќ��F��fy�ͩ�p�����͝Hڻ�޻���m��o��p��p�t� #_�?�U����������<��PU%4�>�����R��^��Q��;���[���X>�3¿R�oV��z��F/,lV6�?�Q�S��J>[_���#�N�(����nJIn��K8��	c��b���ħƉ������/$a��/M#zOҨry+�w�a�4pf��~�7��9!)��8n����S����l�8Ӷ�n6� �\:!-mA��v�T(8��4i9�dBB��QGb�b���e�.�w��kq2�}#B�b��׊�Ȓj����q�&�GB�o�e$�Y�������S[P<�Sš��9�J�����u9�n�⦾�(����<�
e�����gb-2��l'�P�5'�p|�Nڷ���]�c+���wm��
�M�1�u�;�v#�U�ț��%���.\JԦy�݇����5�%#dy�e��F����a/���>�cnǂ���>�q*��
B�,	}3���ϱ�1M9GSegɡPH�[�U�\ew:*}�Ж��� jM~��+�ά���
���P��p�Y��&�"E@>���f���1(�Y>��6Ծ���{�>���)�e�ba]��@��D�����%J�DJ�]Ҩ�����>��4�h�M 
�dL��b�.�����Z wH����;��.٫���5�|J��J�;z�c�d�l6�7g_e��0R*�3B�+(�*Q�"��Ai"s�Z�)�g��C��S��Ak�R�x��x��l�!�U"=���w�5{�����֎%��5�V�(8� ���;�=8�6l#I�f�	�s���B�|>�2. �͍�C/3i��P֒�˹�QiX������zO�cq-�++滘�~��D�)�T�`�J�������%�C� ���,�P�9�l[I�!ې���7p���)�Ȍ�&����`8���Z����n~�� [�_�
�Em��Q��<U)��Q�R��Qr"QZ��h"�Gj��.��
��0=T���h�yB�KTow���~<�QŻ���*�ʋw,�����$�;$�]^J�P�|�s�πds�X��1��>e�(����n��h0���B&�F���煄�z�'zv�k(?H;����w܆+4B��2��	�}W9��6����5�6�8�/-�9%T(%4��B��e�����N�C�^����s�	��$�r�7���R�^CL���.t�8�-�-�\S1&U��ʑ���%��3��M�`���Y]Ht�& RtS?���4�ݽ~��ZO��\c� }�eC+��\~1GŻ� ]�a\�+:9k�v��\(�`���4��֒�d�,bZ�6t�bdK��w�	I�tFW�$=���=15�0X��]/�;�eQB���V���~.:%��k�[F;�Ѥ8�5]���߸�.lt�����t�q"%�CD�CN�>�n�t��晕�`v����������e��ZFq�qpao�j@���?P�%@�S&��Âz3��d���3�ϖ�9�0Z��+\hX�(P����[�h�!��E����6�e�;n�����r��e�� 1�Op%CO�2yT���V{J8�����v�oѮ"�Rb�V�s��_�u��R�"ǋp�C�NST��Ȃ>�n�U顋,9F�%�˨[J��_�_����w� ��ø�~��!��b�����Bh�Z��|<A�@��s���b�~8,_3=Sf,���"�N�f�S����9f�-i�w��8FS.�_�xx��ۆ�.4�	f��6Au���n\%�=��;,TW��EG�L`Iɜ#)�ՂY�����.bȈ�����X����3���`s��ȩ�H�%�����ٳ5I�j_ś�]XkQ�0(+��9FaCN�T�����rm2�
ra9$[�ѺϏ�s���q�z0~N���X��&��a���SʿxBrܴo_N9 �n�	�d��J��o4,�,�17c� ��a ��� �w�D��M�;Ƣ�b��Śk鱯/s�8$_v�`���W?� �%"�/���`8�~+~
���ڤ�Ʋ�/�'"��y3�<����r8�'.�^���k��b���ˢ�~j`��"�K����F-���Y��9DB|>m�d��|#,��sG���<�?+0���)���@V�+�.��
xKV�r����ixmt,����B)���=��/]�itM>/�ɐG�$�7��7(^^}[��{�id�.wPU+�dY���]�i$��/�2r��>A�ӐA(���*��m��tòBN=����	���_�?�E���tDS��.�u=�Z@�/�ѥ�?�g!]l�-/�� ����atx�������?RQ�ߦ�<����A��;�C6�tB@���H�[��~�,D�X�4���_82���s��r-T���*T$_OI�{u^n1_$qw+y��0Ch�O��1��Y�օH�|i(��mA6�]���mif�_���N���f�RY���f���~0{.��;0��c��{c-��
��\k4����2�j�(� ��9>p�p��G4��D[6���0��K#��D�yu���?u@��J�i��V�d�n:v,�;ϫ�������@iL \���(}���Ŕ��;φ��I�s�m⠙jfw->.>����>ϫ���٢��}�>>|�	�- �P��k�4������E�� BIӝ��pZƋ=;���2=$�{��� �ẉi��M�.��Y)9��EZf#�%P�����$Q=�bc͞���\E��G3����e�^��\�c�sF� �ܲW���T@�sK~�~^�e� 4����}���n��݈o81`+� V�_�|Iu2 �ZΈ�ͭ"yI������V"��p'��	�0{��s���].�3�j⋞��y�u~��d�?��&1�		��V���+�j��m+}a��h@P��EV�7Oi��k����村S�-L�5#:��� G�E�2�FY�fl"&���W��V$zG�����u>X�gß+���dd��-q ������ͣ��p���Ķ圜 G���'��c�R�Ԇ\�"܌z�VtLk5�iV���{چTr{���Jg��B�J��o�'�ͺ*�����g���r(��`d�kvV���B
���<��,��ZYRO ��H�ʰ�����|R��}�-[G*b�{J�p"��:tw�
���Au`�L�wз恩z:Ծ�
���'�g�X6f�<�*�q���h>=�]�;��c�弳ʩ����4������`�����W�V���m L�V�sB���p�;ܦw��5�w�mWx٘e�Mߝ��4�H+�~�l�I0���?fC�ܴ�F�S]'��#��ί�gy��D��ߨ�q�g�����Ε���$N	}� �f��X���2p駫�_��Pj���ըO�cI]�����cjm�_���(n���C��'���AǱ��=x�����S�1��k�n��u�5
�k��d��i��ýNJ�,{?�����z�8ıT� �x�!�@���X*��	�lgƏ�9�n���@2X@T&�p+2b�Z��E��E��g�+8�}#�Ȩ@g�l�{̸�<A�����ʹuf
s�t���C�-S��]�W���!`�;���@\�#2	v%J-Q>��0 i7Z�j�R����\҇ќՒ�hO�>|���<��M��c�4B��Xj��	Yu��6���%��J��?���08_`QD���9j+�a��d���
ȀN[.d��OTvљ-`��o��p2X�u8	�^N�ve@�q�i�ri�%�1�H} �hցb/�6u���Rse��p��ć��v�I�E�@1�!G:	(�7zt?�i ��c�=�+/j$	�]����ʖ��gϑ)��n�796v��$b->I4����nGi�il�4N���WU�P�)]H)GW�;���'=K�HӤ9Dc˟յ��C��>����Q뙄IK��)pꑊ3m�����U#ʑ��!҆�(=V<���W,{���1u�#�+W��#ԭ#��T���@�S�s�*`���V�5�keB��{Zԕ�rK�kH�[�*��y{e{e],���p�v�)��v�ϑz�p�����a�a�Ȧ�-�T��RL�~�����C�0��P��`���<�9nd_����-��i|	@��	������{��04��~%(���W�@�m�^5���cq�� α��HF��9�sdtN��^2]q��gN �)_K����.RX�D�%C{����S��4�h+	o`���D �c.X�>lVFM����2�N+~���ч��|J�@���fE�������+����_���Q������s���^��p�������~���{%#���^篒�/u�����OL�T�9�{a��׾}XHs�L�j<[� ��-�"Ɂ$�%�GM�Ź�mp�l%�k\�г+$�.=���sF�o�q�i�����Y��[��
�����TM�����I���6�3m"���"�c&$'	�^d��D��W�R�^R�Q��$�
$�����|>k<����9��T��4Y�E�%����֠�4���.�l�Q چ�	P-���#�����\Zq��ow`8�l� X�$���|�ب@ι��^ތ�Y�\I^=� /)��C���c� �|~����p���+�dԺ��7w�<��x����8��k�␍/�Q9��i�zf�h�U��/�N��� �Ow�o�S�-����?V���:6��S���s9�`"�
��Ȧ�?��V@�\q������rG���l ��b��u�����b����!S{V��X(ן�ѾL����b!j�9�A������0��8r�{�j�Ѥ�NB�N:�$�u�%syv��
>��� �)����JF�ϖ)�!.�:>�8�f���� �}��TwA$(���?����~�]��q�h}�$���q~�T�>A�~ڐV��L����p�UR~�����w�c9�ȭ�'T �cH<t��2����q�d�@Y��2�b�n�ÆV�ъ9d�n���gCOha�AԾ~���t��2{�n¶�F��_%�*�J�o�O��.�I�gOG�	��i!lOc����x#b��A��_TF��E3�-kz�/��}���?�yTä�~_��72F5L�����z�=�J��XD���2�N�<ړ�;�F�0@ˤ��� �&g���!X�n��OT��W�6da��η�ߑ�h��a���ŭ��q�\�ӫy�U	bw�k�Nu�a�75��ٔ�DZ��x�D -}��ҭ�d,����d�Pa���?]]� ����[C>r1��1�
����~0sh�v_������BTۑ��$��|"İ�I�N<�Y�/�o�7���l_���!�#���E\��)��������f
�D��j���!����>�<q�A���uSX�ݦ��#��c��}�xCx)C��6����ዉ�����Ą��Ro� I��t�1w���[F*����������I�`T�
�G�E�t2QXr��,�(���^�L��*��,�z��N�B���k�˒���=����a�R�7u���+���H�N]�oI��Q.��N��
��Qs|��ۛ���J��l�s��g���\�@�'Mu3�h�Ê#�77IYx��&��
�0E
���ZT;��w��?�wS���XXz�:�H�UYNkm(Y+�
��.�3"a�TOd���'�~�۝�������J�u[�1����%/��1n,�v�V�;"n�z��}B��E,)-���u��rҎK2Kd7��R��A���=�x�N��T��8�Z���Ͷ��u[L���-N-*�J�XS0�Mo�C�*�$�+|櫖Y�g�S����]���Ni�r��n������%Z��wӒ��W�/�����#pWb��|�\��������w��Я������B��f'(|u�"S DN�3tz�X�`�����w��y{�o౦�N���Pw��Q�.���*��b��u��Ch}B��$��Bx����l��0c��@9��y;n.%	�OE�>��\���ˑ��S8�AZ:Tuv��p����5��1w�
�����Ƌl�(H�b_7Ҕn������&�;�u�H�V$�E���3�ڇge�rҁ.X��b�֢`k�]u*�@��N8WZ<��Җ�͔�Þ���C�1�I�I�u�OC'���ڼ;}�&�O����ԧ6����W2���/Ɲ�KMW6՚����NCv��@�I���ox:J0�|�`ȹ,fP �E��!a~_W_z���s��,r���w!�A{0�?��G�Г�o��g��Ͽn{���Ճ.LYG㸮�/��ˀ4��rř��-)�F���_�(z-��Z,8�uƮ|�eE5�XG�ɏ�M�K��-��|N�������Ssn��Λ�����e<��0@]����{��A	|�D�J�(�R��$Y���A�Q�N[�"m���󦁓�n� �l5O��VƯ仚��C�:ּ�oM�z�d���͵�Vr���jb�輩�Ob��F��&���%��,���Zi�yC&=b-
��NҝD#f��u���ڇ���k�t�c��N�}��8�Z"��ƚ�5�y�l�C�N���E��|����ޗ����T�����?s^�=;b-����0&�b���l��W�qP���q�&fuL���0egA�)�q�;���Z?���%s]A+/������rq���-U�C�4��&��#9��8����e�(��ۚ�=9n��$q.\�$�����Y�蔃O0��z�u��ތ�:/G��A�t:��������@;��I	�a������ed��YIۥ��{z�ss���ihİ�4E@O�w�AO�\U$"����K��I��M��T������[pF�g%<��>AX'��߉��X��fQ�s�}_MFґt�/-���
��\�e�~^9�����D��Q�����^Av���c�x�g�ΛU�-g?�s�4�3i��p{��r9�cg3ҧ�%�!e� ��Ibs���@�t�����#yL�İ46WR`f����Q~!�>U�@'����J��֒�[��M_��K�����5	��ᤛI�)�Ck�p�B��Q.$����ߚ�fe�&(U�o�������S�4��k���d��;�W���^~�7wt��6�l�K��qYWWX��u���Q�y���;S7x�{��������Y���<�w%熪f��&ߘ��P"���� RL���Q_U�T{F�Q��	�IE��շ'�n�#R�Q��{B4q;x��
��N���Ţ�]�Zh1y40"ֿ6&�]�D�U%.�X{��=m��*�k���Xp�#%f"��d۾�܆d}D Q�;kCGN��H',1������S|�ъb���A�A��*�C��o��\+�d���b�7)O�qJ�Y�|$���O�c�6��T��1C�{����1@x�������M��⋘�!��{5ڣ@��{_m[m��UK�bOTX9D^�@L9�ae9
��K?�O�ʟ�2$���D��	P��ORi+u��m2o�Y4�3��ߌ��ܯ��Q�̼˩m�t�;\脐����w�q��D�����?��8F�WX��{9ac�5[�	%"X#��^Z��BQ�
�7��{������4�]s���7<��+߾%	h�O�ZS[�ݠ�{�c�y�7��ew%6?�3�#�!RR��!�A�ӆ�J�&�>E1�iy~�����g������������5	�z�Z�#��n�`��������UW���Ӧ�|Of;A����{�`��4h87� ����4��"�k�k~���f�� �_���/Ә�E�y��ws��t\�O�Df�W�pmYJ*���T�ާ���83".l��<��v1*co9w��b���^{�9z��[�-��GQr�]��!�bWo��Tɽ�3S��EjhfM�2^$k�Ҽy��|Ж���\�.�ϊ�nN^����o��Κ��a���a"�C�����Ԩ�UΆ�4�5Hl�Z�O�$�-�٧�90�Ȁ*���WXU�E��&�~������_�+d�_i����~�>�toA��Va��#���h�!��{W+Tv`A�q��ih�V��M�A4�PH���O��fb�!Ϟ��).�Po�`����'����QL�"��w��Dc��ֆ�[&�:���V��ڹ�<�/J<ٿ'7�c�'��¾&����=)���`^p4s���<�JF�#l�IY���ÒY��0�N��ݵ*k�(��f&�m��"�m&>TM��\�v`�X�U�������aE�Mȧ��K4f���=Mp�C��.�1�C�����@V����V��_b��g�P> q\Х��`W����a�]��iC1A�wp>�^g�bo�A���"�gV4'TY��7�j;a�ȑ���#�9}��Tm���=A�ϼ,F86ٚ1Ȍ�,��C��=K�2C>�c��b�0Fi����j�3_�!�4C�=U\�Ch{���'{�+E^�e�MO���hh8�^ؤ��X�<r���∅&2b�R��:/C�4����<���c���B9OZ}OI	�)�����4ϋҭ��~�L֮�s?������%�	;6��sg�?X!���s(Z�f���ܢC^�������$ZE0z��3/lF͂�'ē�-�>w)��إ�����`�?���>e6*J��|~j<�9�(�`��3�y�Tż�5	���+�
�Ӝ_˜&�O���<�
<	@�p�����i\������������i���Bb�l�[�渭xk�E?ִX�=Y���ώr��������Z�Hɷ��s���>��?\}u@U�����Cꒂ���E:%�K��A@BJ�J#���tJ#)ҩt���>���?{fwg>S{f��"�]U�d���{J��ّ��ٵ���ϕ���^�a�{č(�H��u,��c�O>�i�Y�����;g���|���5��8y�@�.^r��.���5�y�9���冟Yi*c'֤���b��^,�C
D�J����k���\���:���ƭ:]μ�73oYeR8CkN��s6d�1Wfy��_�y�:d��Sq�}>;(O��eӶ���FQ6+�z�C��Do���r�l�\�~[EJШ��#]�P���<v��-���},QԒ�������?*�W}}N�7� �L��/�k���Ifa���r=�ߐ74]�+��%'���O:SF�v���"��� kƩ!
�<�����.�S�Y��z��&�'+s���/�~b�����W&�N�y���"��&1�t[\� ��{��g	'٦��Û5��ד-�@*�1��px�h5�Yޤ�ў���z+���$s*baR��|�B��<�Y&7.��E��y��WK��_�_��	+��������*���̹"U��m��)%�.y�7�.T��� [��|��@������J��+0�c�>�t�J2&rȳ�K���`mN�O��ҋ�<w��v��\_���J�
Pv����N�t8CZU��J�a����-�L������r:��#�, �˖ok��d t�����VdfSғ�*<f>���?c�"�rC��������{�[�%6��Zh��X��°�2��:�!�喯Z�(��+I�}> S�)k�.2s��L�c�1��ę	R�7���__J&o`&���o��+k�K��r��t&<|Z�����$v��GD���k��qf
:����^8}�U��m��jS���^�f�[@�� , zϙ6��Y�h������ֵ� ��H˖{������-ky)��,|���e^�|�Z_�%��ن}��o�	�XT����{�¨i�b�m�����q���\s?�ٱ�~K��*��1����q��x�Gd"FY�`����	�`��BT�]=F��7�'3����b�p!��b}G��];��m�B޻|/_�˰g�uq�!&%��wC�H���4�oVx�8���tnؐ�yx��y�5,���Y��M�z��Y���0S��T�b�������F?>A�u%���h^���nm~�v����R3���d���{�jp������� �,cQĪ��n��O1�.�E�#����~�6�}wfF����.1�;g&���y<���?����fSج����/V1�U:���.��G:X>������>�^oI���Mx{"�˾���Љ���=u�a�n}�(tALI��!|�w�s��<h�t|�;l]x���ru��<�f$�����ކ넋ll���z�J\�=�T�.����*�J��K�%U���fz��d��~�X�y��u-��g˅�kz�d}�ϭ6���w�s��T>]Rݬ�Ni_yH{������ɿOp=��G�Q�t��ryG[d\�n��>Kyu��,��)r��wl�n\p���J�fi�ތ��XՖ�-r�Đ��`L ���! AeߤБP��l��7��Lfi|�)AX��-Ҷ�g�L�8�ӣ|,�?/C3����Fp�O#P��H�ʢ��}eB���^ � L�L�� ��l��N	��5Nr���=��m"��s�Y7 >�\d�?ʶl�<ߩ�f��֩W3�	���]7�N֦u��&��@�(�Q���;�.�vV3~+���Z�i+� ��5��O��ܘf��bKXr:HI��BY��t����4z���T����˦'i�8�|�
�37aX����羬�R�7�a�}/H'��s�����О�J*�|����該��=�*��/l���I|O��ZQ|�L�ʅ�+��-�~Sv�Q�&g��H��)�}�sr?k�A<"�[��RBZk���>�N[�/	6">�X��Y�+$Z*�WJ*�T(��C�Ƽ���I������՞VgVm�/_��;����7��լ��g�����}�	���:�V��p�%䢟��K���_��'ۛn�bMJ���e]^b*��6�!��'	5\p��3|,-��dZA�S�GWp}�~���U�G�O%�2�����dd�bS�s\!bqqKq�:���m|��T����������-�,�_!�8v�\d��w�d�p��ҀO���D>w��5��
*6�c��օ7�>b#�����.����]n��[�V�m���!u_�`�.�%��#v�u����{��%�����54D!��DF�ؼ������ٝ��Q[�g���RRZs1���f�"��?=�F��VOP~�K8B�\�򎂪FR�ng�^!hSt.^&�p���~�����������Z�t��U7�*v���̾�f#�-����y�u6 �0]�n���K1q�����S���*����N��@>����HK~�������3��mpK���җa?K7��8��_����=�m�k_�A�2������X8��.�)|Wh��*r[�s@N.��V������.�hx��7=��k��G�1�D<V�y,?�f�b7���e���΄1�kv��ջ~�$�興:�P���R!��<�&��A�9Ӻ{�uZ�Vo}�"�;G	�NE��d�Xpy�5��o:�R�	x�wib*�Vp�d���na�V�(�.��j�O�L=d�qpR{��_�E�����*��˨< \��
Eq� �RBW�6��v�2r49E'n��}^/3(��CW���N8���T���#��l�0捍��	�ʬU�6�6��T���zE��fI��kA�sB06�rcB<��I��[���1�;�E���ḍcX�¶	4�8�~��RWy�4�}fJ�ź9��ơ��ݨZC>�h6�Yޟ��Z\?V�}��SǞ����\��~��" ������|��k�:���Ͼ�����w�=k�J�}^�4�NΕ��ϵ��g4�rwRJ�k݈[F۷:�<�WLR!-+X���Ǽzb��	�R}�u�/�9v�{�M	!J��ɦ�{�M�Y&Ɣ�b;A.a2�f�YTe�3сP�_Q�����h�����������=��e�ğp�B���6����L������Ul�3(fB �r�����I�jB�`i��f��C_k�d�^6��ui�=�h�ρ��Ѐ^�-�=��D0wNC!8�`R�bC�I*��� F�Iit�W0O��T���sW��+��'���m"h2ڼ�^o��l����D]�ÈMMpc�1�WDLe��7잌�8�tmF4xZ޴x��i��'��� ��Y-�!�\�^��!��D}�㙹����t�ݧ,e�5��A�=���xl� �R�{�$o��{V�q�,zt*o���7���ڔ�����ªz=�'6E>pDQ�1dS�����s�]N�׺��z!����L`��
�f����4-�)��sO��X5���X�t�VppЈ��7>��U���V��9I������sz�B���B�DS�r`+vm��"OmE����D�2#{hZ���k����TK�	������+Q����H�����x��􏮺/��j;�?�ʘ�b����U7�0W����&J������ZP'����=(������4>>-ٲ..�̘�0�M�&�%�c5F	K������c�̟�tӘ�E{Q³��	_�BS�y<锦��#��5���GgZ�|\��:��Ѻ9%� ���B���h�1���v���*�I��?�i��7y�N.�A����/؞zv<�)�<3a�f!n��syM6�͞�FK	�I�_rS�'N&�1�a0��OI�9��Ӆ����ヺjĿP��� �G�����|��]�)"�)Ȍ�E[���]�	_J�&H�\��D[?D��TA~�[F96���}��"M$��(n�dNqx�Q�i����+qK��W��h�܃��c�Vԍ[$�A��0�z3?p�\?�Zk�v5(�0%��6���U:i����&e�#� y�Ρ��D'WF��fI�!eb�����(����++�W+�ѼQ�������D���֓���p�cx�y65l w��Rk��f�L����]���?�M��K�E `5s%Ϗ��x+���E�&���~7�}Z�E���A���Fl_^�.V��8�)�^��Gɧ����W��&J�-YcL)A��=>�=b�������λ�K���oR�c�M46c�8�+!'�N���N��r����0Q�BS&���v_kF�E�;HBIFS�a�^���n���/��4���H��	qs]h�h���o�]����d@t������_�6N���C�G\���#i��H�Ӆ��,o����ʠ�E�t���G��Ե���� Q��Ս���� �N�ۍ�˦��qm���V$?��:�:gAE��6x�
?��}�7���ړHD�t��a��)�Ay�5�ݻPlp�����.�N�)0�|�2��y�%�i(��� 'ʕ��]y<F�2y:��j��Siʇkw�ǌ��a��Mw]Q>��$E-L�A�-CK��ZN&��$e��?G~~F!r�q�^�T�-~���̎�?07�`@�O,�L;H�6���:{�	�O�F�]Q2dV>��`�:����JWM�7S��*�U�N���`�{�?dG�ąl��b8t�ʭ`�)�tvZY��&�£]�S{/����U=�y�-�j}�׽���3A*�BN~9�)?w��ـ42���"9���.�8.n��ۖ^ XI3�\$���T��LΙ��*L��()v���r \�+�II��?��<�����;�-֠����pb֚��%6� ��CV#� �~�%f���X�b�{�����[������agp���D%�']�$x������K upϦ@Cv���u���h�:(���#�y�'7�|�XOZn�T����-��A�3�t��U�6۳��#Hp�o�&��(|�@��ӆ>sů��� �^�yZmJ�����k�$� Q�zt�g�:Q���=�_�pĦH��h^Bj�쪢J S�����{eb����S�i���*����i$x��Ł�Mz��k�cL����b���U���sj8����t*���%�`�>[�QOxĎohkK��3ڡ��yD���=bv1LF1���W�O9û�n"0.	�z)�c�U�u��v�-ı�����#~�BC�֛��7q�p�KRgt����-���G<-~WG��-:�oh��e�|��u�*{M"��qI��~V�3ad�iNDH�ɞd�Q�]}@�)a0��UI:q�;��9\�!5v��� �ֽ!ܕht`�388]�%�ʶ��@\|��e������(��!�����5H������X0�ڂ�%d�g��BvKt��|w���'�7YV7&Q���o�u{�I��Қ�@�!\;�B�Wkn54���ar���L^5=�t������C�l�9_CE�O��-1�ѪK��K�ڱ�T��n�]�z3�����*�~����v���PrE��e#�2�5.}R�Mm-���}_AaZ���.Y��������Y�Ve��SD��X�qQ�#���P�ј"~�?>F���^ #r�z��9�e��I0kYb'�:�7�)�dsE�w7&Į�,kp���s2��T��ŗ��'6ş��cU~.�"��I�S�b�**SB��G�Lt$H�;]���B�
Bˉ��v�>�r������R�iMB����۷ 	ׯ�2��t�F *"�I�!ܺ<�K� �"V� |
2�$��� �w�p��%�R���CMv�����J"jE�b�ď�?G1'�B�G{�0�G��#���*K��"�?���?T��6�?�M8�UH/~��59���57��Or?k��3>O6L���D���M�D�(u�(��:��fr�K:�!��V��8��R�G�]+,��i��5�3&�0Pp���<:u�1���+ }��|~y�� �j>kx�ӛ������U0���ЊɄ��&���al\�4ݰ��CƁlY�0K�����췳U��~��
���X�s�*0K�?��0�v��/M�d8��p�9�l��cjj��;��'H��ɾR#�Bh<,n�ҙ91y���s�U"���Z����GD��r��2��c�vSW���)�ΊD��:{�}c�R��F�����?�K�+�(rb�N!��a������3:[�LӾ^Ub���2訖=Qq�s�_���ya�k�N�i�/�<�?FQ�џX�N���
i�^�co����nyGA\�+#�C��K�F�7���gl�dA���cTAl�n��~5�BzB��6�"����1���ZJ�Q�V����L/�,T��ߤ_?�-�O�
�{��c�i*�\��Prv[EB�a{�ߚ!Pۭbq~�\q���w�B%�����8�A���fh��Vט��RF��Y��H��f�;�)"0f���栢������p��2�P�$�?7���C�o`@���&�B6]�<@Kc�xfI�x?�ц}}1�9U,	�$�<�u���u:>-.�L��ᣞ��|M:��1n8ls�b�<��-��R|����x����%�Jan��
�%Ww6��}�ѕ'��9���+Y�q~�:1'7���y�CH�.�`"�\�1��&`Ȩǣ*Ӻ����9���ݨ9Z�z�Q7@$�F�x����w҃��y��#��Q-�m�u~{��A�r�P�����%R��O@uafU{x|�q�5,�wqG��2l(����{/�	W^p����0l���}�Ml���e���9�5�0���X����t��]-�#z�4z�mw�L`;"w�לY[��Y� �;ZZ:%��J3[%	�����6ƕȊs�g.ފ��R;9/]t'���6�b����k�W�)�%A�}9n̃o�?P|Bi�Ơ������V�bT�-�c��WW��*����6t��3�o��IԨ��,3	嵝v�9�Y�^�^T�5�%;��Z��:��cR+p��YC2��)"R�%0�+>d�Lڥ*N&�H���
�؋�F�o��H�j+��<��7�i�͇�Ryq��,�T5������P��nIF	�_�!T�*�(U��n_,�ۥ�F�Pn(mC� �v���w�f�m�U�1��柋a�֩`�i7Ó�w^�}��=�a�i4��N/����k����!.=O`:HS����dE���m���F�0�&�Z=^w��y�����/rZ��(�7Z�M��=��Q�!ܟ��F�#�;<����gL���d�*�"�z#�g���)��E�^��|z��^�^�b��Q^̱P.�����J�ʋ���}ܻ�8��}�8��Ti�iG.����9<���Fpli����3X?���FY�aB:�����rz���!��lq��C�*e�f����e��Z�^�Xϴx11:�"$Sz�'� n��>O�*Hd��2l���<�q�<Ú+0G1RT{�-㋶z��EW-{������/Ԯ��.���blA�q{�K���S�$Ƀ�ϫu�  و�[m�io��\���Ĵ$��9��Mւ�`�$��XzM�mu���*����P�j�Y�aeBXX��b���yx�z�%%jY.���r��c�?�#�]�����-B �%�E�՗�T�<��Jxgk�
�M�L����SU�jܾ�Z� �������"�������9��4GSB7ߜA;��9�eͨ�BW˛��W92K��O��F�<���Y���cz|��?�$���Î�ý���c�]�(��i�A���}¢/a;9?藨հK��f.׸%j���3�}�F��~�� �<K�8%�B��'�7A�>��Ԥ��;��St\0wC.W��#��K�W�E��zއ�8��REq.��A�c�	���-��L<��xJ6H��]ۮU3TML�V{ź����3��f��K�0�ĔG���'���[.lR _L `���9��\�j�I��(����ӭ4)t���$q�@�a�	� ���n&��Њ~D�V��ݼ�v��e���^�e5~ݳ�~=�#t�	A�]�=	3���Cq�ى�w��7�ʻz�xD{�	��WG���nF�)F���G�L�7��\E]�p�,wG~����WL�g���ೋh"tI���N|��k���Cn��a15�P�2߰ Lτ����)�s���¼vߤ	�f7�7��+��1Y�Z˾V��𲲔���_����E��gS��P�7�l$(�Qq�|�O����� �����j`cљ�'+LO
�0�����i�8�h�sٽZ���S������|�:˧�A	��Db��hy㮅��rݗ��aj=�?�ԙ/��+IA����'6T7 i��qO�6{-�>�R�~7)�0���0��o,1��B�������\�!���#Xb��P���?Z�m���>�r��a�D?�B��x���I[1���3V�I̱�����L�&CW����8&B pW$P�r����&l�����1�)\����ѽ#!r��)�A�i�L4f���S<�MV��>ۆ}ht�V��U��	��!��zy���kS�nt�j{廰����i��a�RD[4� �'�kh�	{��Ź�/�!ʢ�<�5^��D.���@�Q��o�r��w9,�k2�\<�=�/�vIΡ�8��9��%*�������v�o�[���w�]��s��=�a_�N�G��2 ������9��.��f��S��紦��os*�>[L/�߸#��.���� ɠwݪ�A�h�g4�( ��G��
�9���I�A=�� ���\,��޲ �PV�|��D��d�_����|B�{]ks�ԟ�݄�L'�O��4�8���G�0F��zs�1��J�5"�!����҂<�_�>O+5[ǘ���{;��-�0��-"t��VDƈ��V�8,�vT��y�Df���-��z�M���K�/��k�@_����+~�|� ��[\�M��K��#F���c����j͹��1X�q_�k<�<R���%��(�&�����6�]��<+�*e�<eok�w�;��߼�Z&�H�ؤ������nW�o��KW��ܿ�j��Ĩ���@�J�i7��	簃+J�eל+�4��2��<�,�6�PYqb�1��P���	�pkB��ư��Ⱥ	k
v![���������	��NB�ѐ�ׂ�Qx�_ y�e�?H,��[s- �+l]Fc�q���/��s��(q����"��3��Q�/[t��Js��O��o~�>;�*�#}��pn�s������`�r�1܍��~	�S�������V���dO~Ò� )g�v�<��wm�[}Qv����=�E���-(��?�Ru�Xˋs~[:)u4��K"���2C�F��\��s�~��/�����	���A4��3?����8�Kwx���YN/�kl�i4Y��^p��;ia�ϥ_ �	�jҠ�G9�S�+��$e��!��۵1�h����W�C�/�&/L�͖�ʉf���q��{J0>DO�\�!+�% M����jZe���0g�`O�41��ym�T*x�kL��^��GL�s_Ȟ�������0D���^x��xk��g��#�Ñ���}cI��YN^�o2yn�E@�"K���������MM��-Od�C�A� "d�|W}�����-�W*�Q�r�� �<��.��]���Q�3�T�]au�zu��1�?s�x��0Ϳ��Lcb2X��)�gX�U�0s ~13R4�1�s��+ZĦm�e9���,�/�}��=mN<���#l*ڼI�,+�M�ٔ�h�4��g,Ѥ�5��}�y�G�i�qO���b�,���h���]r��. Sj�s3p�p/�Н�-۾{����m��7�8^������t,�oZ�e��kYP���R&6���n��9S�"��02
L�N�����kOi�e��J�U?Ȧ)��<��(
$)]�`��1D{Y,���pN�r�&lO��� �@(Ya�S'�*��1-�����|]@����=n6�riK�Ș�ڬvi+�D�m�҇�q)��&#�jvq�M�!�CN+�)bP+eN��fR���=��c�
<Ǚ����*���Grw��7��D�ќ�ww�z�P�пy!�{ӸM����*5TwH�*��iZ�#w;k�6}~'Ih�쏀�<r@NRfD�<;;!�_����?7�j�c�7����F��yۓ��/+xT�c�o�j����kZֆ�J
�k�_q��l�v=��G��͘m8`��������c�+��f7f��V=�˭E��FT�.��k��څ0�w��,����ߦ)������['�?�RV$��C��y�E�hR��h�8�$�m$�޳��a��1d�z�E�;�9j����D��H \U��m�{���v�G�����I��H";� �H�u&#7�v;�`g�ny�?��$��}��2:M�!������-�x0��HD��*/k�2�2������߻���F�h���M��
tJ0n$�W���B��w���D2�o��ҮF��?����Գ}\�\��^�8����QQ��;!��es��;��24b��XY��9�ϟ�9U';��� 8(�O���>���!��-�+:�m;a�W���\�$������oDRRgm=7:�]� ��*+a^5�Ad���IV�	�D�Jpt,��K(mԞM�^�ɂ�����}�(g��bnL3��g.��7�
������t�y�����CaV.T A�o䒼��T�a�~��:�Dl��%�Ǵ~�w�éc����C���x'�"�]�{m��f""O�
d]#�5\
�8��5�\\�+%=�y�m�fՇ[�[d����^2�X�tzr��S�w^�c�	����d,Ee>�lb���@?�|iD���>������W�O�E�b��-�yVA����}IJ��[��mz�����u=�WWNc���󵑔<�ئ�왧�Cz�A������zgU.,v�V�D���'�#�f��	E��h!5	ހ丩���C��XB����hd4�J?�����a�;'R�%iφJ���zB��-C3�M�p�����1X�9�e!H��v1���8��q����|Ko,�4����6ػ�����e�H��m �'��17�nCA\<�ҧ�����5~^3O��s]t�].��
nn�n��}U`IL�6=C?a�ᅘNLG�E��d0d`kDl�WE?��@�@�JO#꽵�ϱb`�~�M	�Pχ&�{�x��I��V
>�;GVn/�FD	LˠV^�v�q*"�߬P��R_8#٥\wiX�:;K�9=)����z���B�C��c�C���D�P~maΧ�Uy�_� ��K��Q8�j�r�����wB�,������X>�N�]�MLZ}�< �<�P����
J�>I��B�t�&[��%3����V��Nqѽ/��y2[���K���%��H��w[�'ٮ�H'W�jh����ﾼ����SUCcP�����m�W��hׅj��_�� q/�l=\�^�[�O��9!�{V�<=}���x9�Y&���p�>ۣ[�/2Fk֢^E�Э����Ah��Y@�L�O�e�t=�;��*����~\�$��C�y����Vxfc=U 5�~�� ���E;K��^������~�|ǧB��V����&�|�N����qτ�<w�̻���oj ?[o��T��X�=�G�ظ�S4��}6t����yL*j��a�OHl��|#8}��J����a#���#�lW��TK@��	*�f_�y��`����!ˋ"�h���r��Y��-��;$L�|g�>�f�t��q��Y.��ќe��5}�%�N�� -_�h�u!^��ׂ)˭��I>Y�7<�c}��|b�$!�8�(�*U��y�d�U,t��(ܣy1�q��9`�G��r�;s�����6��f���^�,a֐��k>�s'5)�n����\�]Dޟ!!ҩ����$�|���O0=��)[2��H�g	�����<t���@�Q�"*΀S!Ԥ�3�o�.�;W�F��#T�ue>AZ3%lW}�,K��t藦=���_��881ҡ�G;~D5q� ���?�職���Dy���Sk����Ib-�K45�d՟��_31i�?�;O<"�m����6a�Ju��e ���3Q��@`ɾ�}��M^��f�/�iw/2~����%��͌3��z���>vj�H�ʜcVw�g�S	�vu���V�&*q�����?J�K��CVbS3�Z�D�a�,#N�tj� �n{m9��g��������*��E��dr��y^��L���kWt���A0�/�G������m2�~��U����6*	\���&�#�7F3PB���L7G��O���q�~z0���S��>0������.5� �<|ztA?�Y��o	Ջ.��ݯ�䟤�5�\/�����ݿ��o�!�����=��_:W���վ�*�'��躿BT��j�k�'v�����kɲH���wF��y�$b��	%��ӄϕ�m.��h�������X ��Ϣ�Urg�0��w���L�g����g�P1�ޭM))�����y���m#���)�8w��ݳ��'}#fx/Sz�{�jba�BP�a5`K�2� �ˉ�\]�oa�C?:4��dYp�{�F�A��z��� *�c��}R�3l��u����"����Og���޹�{�*-K��~��^��3T�A%����Q]�7��2#���|�1\ؑ���O�u���&MK��1C̥]/Gp��Vio����zy�6Ņ���b�!�ý=Z���Q������=��N��%��"&^��X��w,)9��uF�R�T��C>��,|ks|�$e��Fw�CC$!i����ы��1;���f�ŧ_�����^����`'�����X.;��mh���TU���f�S��)���+�ǚqٓI���6|�Mk�)tGбx^��CP�#�nTҽu���'��&��4v�v�N�v��Ad�!��ax�ad�ad������D�m���*�A�/�נz)J�'�'��sf"��$�m���a@@<Jd�I���݋���^�P�}�ܳ�?�����/:m�;w	�m	;?��!���=Z�2JT�k�L_��K��;j��St�Y������mtL�fz�h��8I��N����OM����2�M�)��"���'���vH9�d�y+�7	��c_�G6q���.���3���fa$�7�Q�M�-���SZ��Ew�����jO�x�$Nb=(���?��,����ZΩ�'˂O"<�Y5�*cC(��mf�:�f�z9�Eve��L�W%����_�M&�6�U�fX�E��ms���k�[^�z(���u3��.��~��.�ɨ�!��������r�M+,V��7����O�#���o�CQo�z&4D��?y�t���b7\	���c��;�ja]c�T% !9
�eG*���`#o���W�{/��f�4�lm�*��-��������2D���*��]��y �g�a��R�b��Oc�|�_&�^K������ �KF$�iF}�јA�����Un#��u�"�&��ήV��'�O#a��'I��k��
�ۼR�c(E}�9�[n�~��m��ӺL5�,��+� P,�M���`����H�R�07>�8��x��Ѹ�� ��,̗B��oo�M|���j eiK𡹃���	�_u���[�u�>م}���I�[6��n��|��A�R��*2~�����?l����s��O��!��>�o�+uh�"�(�@S�Q�ͅ��ᓺ�K�1�#���������QB�$�J�����W��o�7�����no6���{����}���{�5h����d��4k�x�u����Hh��Px�id,(�i��?�i;)��9��A\v)����,7\*���S���<����)�9�����zv����[�5¸�ƮgɕG1�([��)W�^�"D1�%<�&����_��|B�Tu-���zBx���������T,8���V���C���,�8|w�TdL�D�5"�$��Z�*�B�z�&���.�w�Y��9#O(Aq�'�qf�e]�;���W�]:�	��?��#��_b��1Sʨ�Js�"�N��b����
aW����t��tw���r�'2��3_���=�ye�M�&����Q,C
=kyR�]|�u���ݢ�j�����<B�ǡ����lVua������5Y;<�EPC��πn��A��?��.nk��P_�a*�!��R?����
���0\cŷ��Y�5/lj�j�;�P�@���/���Z��&d����pꮟ����?}~KT��C�_}�w��lƝ�gV�J�h�{��r��نP1��p�Gq���/�V#%`$�`��겔���ߴ��*�ɻF�d�󳍍���u�2082��?\�"-S/�j�չ�+�t�ޥo�4\������j�w���
O�������
d,"�D*���3�2Ǟh���P�c��H��hڦ�ӈ�����!���v/�v�B߳r�(_��!�'���N��!����҂����i]V���ݛ��؈��Ki��>!�� ����J`��F��n�7�@��R]N�6]��a`1���BV"�T���U7���(QϽ\�e+� ��ِ�ֲ#��~�C�?���?�[�=���a��%")��1(qz�.��x	1zny�?o��}V+��K\M>k�h+V�I����pwW御�4���Ӣ�;1�
R�F�.X�vj����8�Y����㓄�b����������F�0��<�'��_+�Nw��K�oh�i�]~���;;��P;Y�n(^�9V�h��(�g���n^��~\��T}����7��wд�k�m�(��E\g��y��ܴvU�WI����/�<�<W����/�	��ӣ�����T�Ry8g0�G�'4ӟ���PQ�"~�+�OUz��hsC��� AU�/u�ڸu����F�*��������gO���o��C֜8|�*���T#~,(*�2u麇���8I�	0ή�*܈~]���dxg�(�TV��Gl���� ���u��fJ����@h������M���*Ù\<��A'�T����$/]Y�`�]*4��['�j�2:�>�z��ujp_����tf�gJ�p�3�������o�$��r4�ɨ a)���R���k�U���4�wު>��"n��-�~	V��S�5�{9�m�S��~n�����(����ȠqaIl�i!x�A|��>��Rpk'�� ��b��y�KI�Ͱ;�^�ji�g�9��}C�1?�IS����+�60@�ʖ:�(����rx1zӾ!�^(�w��ΧԸ��b��S@�pr����)�t�� K������3�Ԭz;o�OI'�{�3���妍�
�ӓ8CK��3�u>cʔ�s7:W��.ۯ4g)���%b�N6k��K��{N�������d~E��{��Ln:=%d��8[1=
K�ME����;	�_�Ǹh�ե��OP���'��A���ꦲ���4И��ث�O�>�a��0y_�d���0�e��9���!��}!�ST�/f�RU ��X�'�ͧ{J��/AG*�~�ŕ��!̲ٴ�L��V.,�N����`���� ���P���X��x�N�A�M�J���'��i_��}%��C���D��{Q���d��K��/Z���%؟�M��yex��5���.a��߲�~��$��6
������.��KS�G^��W�?�K�>�~���=��ۑ��a,�r����~2{���	_X�0�P��NA����	�1��8�O�g�4�_p�zJ��Ǔ�������Ԭ\��i?�bZ��S���K\E��U�n�L�擈�����x��=�H�M��\m�~���@~`��Õ�g�i�_�"�V�L�����r��m�����=)v�����H�q;Ӭ	�~
>�=A��57Τ����:�'o�1HU�-< Z%��z���%۾�Й�- BX�QY�їP/�K%�gj���O �I�`���g9�` R�x��A��"�L��{�	M��0��Tx����s΄=.Q�T+�f��P������F��w��ĶRZ��n>
Ǜ�G$<%�
��U?J����bT����(�isM��o��~��}���*��4L&� ��)f��#$/�]�H�s�}1���ӓ��y�9�x��6y�_5{D��'c�!�;�mb����nɖ����`��M���rM�]L�����<(Ȁ��1���������~����K�b��M��V��)���L�ȔDI�xG,+��8��>�N��4:���^I�Zo�G���T�Q\[p�5Ӟ|��>�����<)H�1h�?��t�P���^�V�)>>38�/�<���WV�z��"�V���ͫ�E�*y�xʀ3`?\��r�	?�#���ؘ�|�&�ql�0_��ȳ�)�͐3�=��\=�����f������'�5r�8�p*e��&���WM&3���n4�ƥ��=��EU]���:���i�3�Iy� �Z��7F�gH�	؏+��2�̾cbl�e?�%�hu�6���rA���6�5��."ؠ�/n�\���ٳ����y���ޏ~�e��m�f8^�����%W�uTI�
�2��|��d�W�7���Q#�B����W�vӉ����9��--�)�։ w�٦ݥ|�����&��S��*
�<r��4���,ɣ�+`J�7�	L�"��>�^�����r>ǵ.[�X���Ѝ�D��XJ��k4�Mo���˓��C�G��� ���վs���>맜��Ǎ��x�ݞ�gyx�G�<�;�k�>$fؗ���-�	>��G�������c��Qн��x�hx�n���z�[���祵?}4st"Gi^ƿ����>�Ęn�!<*�i���ѱ4�D����G]�EIJ�7�-���k�`��^�U�K#�t�
J�4J� (�݈ HHI(")��]C�
�%�3�0���=#���_n}����ٱ�Z�X�\/lY(��7�O�|�FZA.;�w��$��e�QwV�"�� ڑ����F'hL��u�TWU�{�s�+��qG-����t�g/AަJ�	�T|O��g:���Ay�,)�(�����ܿ���
HF୽��_E��p���R�j���O_R�OT���g��>���1g���ݜ�9�\�I�� �e�������-P5�!����s���R1�c{&�r2:M*�������2��h�����C~�?��&Z7��E�m��)��>>	OoU7���Fg��*U�/|���yn?	r���G ���c���/�Xј��zU�Ϭ�2��a]Ef��F^@��W��is�W��Miz�s+��lB�.����cSF�z%=n���CR�An�����[��nug����]X��F��dy�F3|����1�.B���1j�������nW�%Ⱦ�iZ�9�y��>�^_A���[������דe��V]H��X�t|��ZE��Kq�dp������iⅦ�,�)�!S�U��@�5��8�F�CT�m�r��,���,��?�b�gb�ˎ�.)D݃�l�_O�Y	��%WO�1�\��BD������f֊�Ņ�/�e���Ҵf +��O�4����k~�:D����Cʫ����W)�\*EU��\��D�j�&|�]���KMy�͔��m�{�1*��˗�e$��;]�qmU�alg3Uݱ��,~A��5�vp�����Q�e+_#�pc,�/Z5������5J}[M�<��y��x�OF��\6U(�:����E.�')VV{�K������M�S ��iva���!�o"G��@��YF��O\o��������nq!���P̐ʕ.��\4+ox-��(B�~;��˄�}` \U[����k�TEI��y��ˀ|������77�#pdJ'�Dͤx���K��ROFCYdFy��!c�I����\�PI�:A,bqٌ�ht]eM�'ϭq]I��٩\�q�Gj;\�՞��Jѻ�=?�"��+�����v�"���~yC���U G��=dK��.2�����1B��~D��{�U���'����,#!3�Ճ*�����rt�\Ԇ`ݻ� Zm#�@R�
�0[�_�?��J�.��Qj��e����A�:9(��db��]�u�<�-}iyp����&6�?b��YM�: +��G���wD/b�r�Ju�s~sͷ
�'�2oq���L�5��e��L}��F���8d������q?����.�#�����6�������Mu۹���_�>�f;��h} '5�y�*��*����������H��_������n��
����lw�w��7��	3��6��i}��k�2O�3e�u���N�����:����"m�vI ��Nu�7����w�s�L���)��C�V�PB��[^yr)˗X��zO�&Ȍ,��U,����p�z=��չ��NÞp�rd�i`-S9����^Ď���r�aVS�!s5��4�����,~����i��wK�eR`� ]���\��ت�^y�L�E�õ������ �z=-�z\��aP��iH�� �\�U�1���ׂ������S��S&��531��ĕ9���ޟ������z"�2���Mv���U��G���Ow�~U�Bۑ���4K��D�/|�hj�]������g���a�����/���a�}{�O[OI��g-��s{T���g�nʴ�y�Z��^�&:��ͱ�Q���+c���[z=!mw�𛿱1�-����T���&+�,"F�t�3���Z2odo4�j��F��ӄ�XxD�����p��͂�i�Wp��W��� �F6^)����c��w���	��$@��}�1(3��7Yf@m��trr��ڲO�+�/��ZrOW��H�r��?][��j��+;�q�y����g�E/saG����/��_L}�Q�Cit��c���S��T�����`!�4ѽ��}�l-���u�Y�pB���]8=��>|��a��ͥ����}��gH��1A�W��A,vֆGG ��<˞��l��6���т.�+��yջ���w�[� h�/�U����⫧sn�N�M�ʛ6R�ͻ93���߮H��z��_̿�2Jس]��`��s<d�sW��3������9Y��ֹ�M9�����L�ҋ�x��� �C���γ��]�����I���9��R���j�@ʗ�Fgǃ�J
33}��s�z
�����k��8�z?g777L�455O�p�3���"��I��)E���k��F���F�L !�`��@/�L��WUUV8�z���8�C�����#� ������$�Ȅ�@Y8�7�k�$��dS��p��[ �}���L��:�U@���%�� \�OL���Y-E�����\�ę�,��:�� H����7jr}�@�]��ۇ��>��!���&��f?]3.@+m�n-3�,���-�4\�[���B���&U�Lc`��"A��h'��JS�SE=�y��'A�:�T�?������~������s�X���>����Ʈg[�E48�Z��`���ÍWq��H��W�����`���x��V˕J�}�N�9�Mo�	��%Gx��)�ռ��(��3+`O��Ҫ���]M�Ϣ~��Z}�y�<&p5������/fT�0��ߣ�|��99�z\N����X�X�u�I�gx��2���_����z���]��8��<<c�*_��5���թ�`,�� ��~B��Y i+��[�b����@������}!�S�0=��h��D�)�0���׎��A�3|��SԵE~�<��_K<^�D^��`�����C��
���$;�fϚµ����}ĽN���K�.��g�$���6��V���q���s���t0�W��Q��g^�4�&��a���r���3��i��ڴ|�1��x"�64^X���m��ϐ&>`�j�=��x����jLC�WCz��Q�D�v1�-���ũ�kG���wvvN�:� � CZ ���fE�X��|#�3��X<�k[=�����k�ͧ_�D\�����?O��x8/�JN��0�N~�;�ڝ��[��ɣ��Eq��)-������8f��<@p�| H\QQ�@J`����@�l@�>	-o�� 1�i�H{��4�X�;��UYt��x퇀Q�K�9(6��������q�����;H�L��*�Xz��LMna!WsK��yFX�<6?L���E�����2I��T�!�@�y`d
T��:ո��kl��p)dɥ��M{/��f��[Vѓ��Ǆ�����jhX틭��~���y�~�+�T_,5/>V
3p�Ó�����rw3�z���m~Y"k��֝gg?��{A�k���wW'QF��!���W�+ͻ��Nm���ߺ'Ҍ~��)#Ԅ�52��~0��R����Ih{��X������x:�ڲt媤$�:�����PB�x+��KN��
Rͫl�.V2�GL���|´�9w�YA�m��@ʭ�D�����a�?\�[�2���?o$�5��l�>�)0n3��h?���:��.��o�(m��hw�)��P�G	@��~��^f/K&��8oc�b��=��V6F^� A��^���1 
@�[�/�uD��|���G&���g��K==����� oaa`�oS���8�Rt��?HO����3s�Jmߤ�`a&`ΐ159���mx����lfB�fMol���f�L�3��:�����:##��j��L3�O�3��TJ��G q��1eg�6��(�����t�K)���{8&Wmm�_/@�;D
��J{9��dq���ބ�[������v����?a�8n�qo+u�M��T�Bn�y ��o������un.Մ�5..�S-�jF=$止[|ǔKݻ�7:�i�5�@����Mc������������7H�O+�*��Y��ζn��:;O4�&�$�P弘PŢ�H^e5y.��(����g��s�,O�&m�pn�5�,.���s�3n���J�%[��R�2���kz~�شl�8��Ē��h֦�v��Cֺ���~�Z���KRc���N��Q�0�u�������v�U��^H�e-n�	�oxJ���^sm��rrTd����M�g���6Y�W��!��5c�����H:
8�q�b̈�3�1�<i�_�mEf[�-n�O����ɹ��f��� غ���y�
�A�*�����Z���H8�R�҆4`�3�v+!�8�M�|9���,�"P�W�Ld�ᒕk�\�10hZ21�r�X�)��/rq
|����h˰ޯ�´B�m/�����"�)���.�KY�;���G,#�N��V}wd�
����~ʂȝW�_�FX��G9ۿ{�I�RGD�Q�A���X_�r�$�̥ԫlJY����|�r|p�Q?�hU��u��C�i\򳑫��*�L�!?h�U\�O���m,,sm��q���J��E����ҾK��Its�#����lW/��1�8�������?P�y���M�2]-��s�nӬ7���>�̽W�gNa�/O9���m]ʠ����������%ޤ��z�;� �ޅ��Y��v�+�G�I[
<�b19(ʴ�nwC�m�R�c�'C�;D#���3J��B�cY|��o�ʋS��f��ϛ������3y-�OieE>��L$�юz~�{aO�*h^���-�r8�+K��0g\g�|A ��/�� ��K7�� � �>���mh�b���� ����x.��E#�k�>CR��t0ا��Sʮ�`F'q�-��?El��R[�>��]�*��΍~�d�[�	C��x"B>���,�����6��H
GI�5���O��}*~���<�q���#�[�,9q�r�K�nd|������@�����K]?l%���R�Z�*'�*�^f=�����5���)Y^����?�\k��߷��T9��q���P�:O߂��d���"9s��?)Z�~B�Uvϟ�N�6��	�&��2�w���v�r�/��*�9�X#�&r=Th.l��8D�,]�d���y6X�֢�Gu��T�ȁ�H� ��ʯ�p�"���)�Y�^�j�^�.j���st��o�	De���S�������4�mVr�.�B4������N.�=�Uu�ߛ�����k�`�6��? ��uD�P�j���B�em��.�T�3b�ghIRjv��n00�
��wH#��i��s �Q�j?k��%�V�(�����#Qtm��ǝE�W-�4��JETĎ�ϼ���Vg�Y1ί_G@����Yml#^9e�3oT�c�
2�Ł,�����J;9�3�hE�] 9wO�~���f�*s�b������<�W�����ͦ���~��

�d5V�E�iv�hme%�	fP�"pe�|��gqŶu�E���>��Q]E�$����Gn��BaV��� ��R�6���ry"b�%�yl �P�t�-/sD�:;۽"7�ZX����Yj�k1�����4*�T"M��P�wZ� K�b�\�j]��!aΈ�ð�Ŕ�*��a?������~<<_rdPN���K+d��"X���Om��-��?9���ӹǛ%(We��9;Q/����DR^�Ŗo�*�i}5�U����|��H��o~�P>��5r��j���X�`�gzX�X����{?�����#���w�J���h������z�c��}�n�{\s�B�t&�Cs:����j�3�'i���)dA�o|�0����GDaM�'�>R���l�M��̉�[^�j��8#M:9�T�����P�Dٝ�>����#����{�!0?�bv:z���(��3p���X�kR��E��ww0w���G0ݠ���z?c�|냜q1�h 4�66T���#Ng�A��l	�u�ϒ���>��`䂆/'�%����t�k�����3�=�ޅd�=��4׸>���6kP��
��}�y�n�g�g���0w�0�{�}�I
�����XX[J��J|i�c�=�SI�O�ђD����^��k$`o%i���'�<�(*-_W��K��� y��aE�������9�?'[��NF�$�A�J��*eB� K��x%�>�y���msP|:yǁ��૥��f)1��>�~�c�i�^�ت&���	ϫg�Az)�v-�@��T�Ydz���<C� IFW�[��䠵R�%���\����i��߭I�/7a��PH|����]���g;J��T6�t�O�n'��"��/E����>�Xճ%'r�i|7�|��_Y4���PT�%nc��
���S>,�C챩bM�L������@Õ}�eM�/�i>��%�$ �3}�#��o�m$5�����<9��9ڱΞ���S��M��^��]����*,%i��vs ���~g,  9�����f�b�b	{�٫�"�E,b����[�R� :U�ٺ�疯o�9�H�����N�S!�T�w�����W���>&����w|��Sd��Ծ8��Mc��l-
��
� �%2�WY�ygb�T#*�0��l�{8�G`��H̑���3$����
`��2�<���z*�+� 䂓 P��ް/?��btJ2�	������.�"�ڀ�bҬ(��4�m��F��d3�Cy?�j�NF�f��O��Q-ЛZ�}B�#��L���޼
�5�i#n}�҆�:�CښPh���ȣ�L�|\��:��(�Jv�[Z���g��v��)c:xiy�,>��<6�W�P�$Gp�B�(Uu���/�ǧ�XOe׸�af�O��6������k.
��}
Ծa�\=�pL*�����=1W:������$D�ʣ/lxr��nk�����'�yhs/O
]�[��ޭȤ�E�Pw��i�}�/�1��_�0��0�U>{��@V�8�l:�s��M��?<���H��B'w��&3��HĢ�w:�m2�t��u����L�Ibn��3[�gKy�����:9H�%@� �Mo�/9�s�L-Q��ܙ�T�J�=J���8�}�}��T�����'_H�Iu�RB�����}>4� ���D+pG'�2�	��yR� hQ�������x�g�I��#؈j�` o�����y�4�,w��������Uin��� �1{����"��/��%�@f��|�_�N�҃�;��g��|�G>�8>���C,�����7����\�S�	��Qi^v�[�ۯ|��lu��,��n'N��T����f��f���_�SaIĢG��ʖܑ�I��#�������SG��^�]r?��|��}�{�
]�����s�z��%(��/Z�ο�mݴl�JӮ��y,BZM�|�����k�����O~Y�}�ĥ|���E���ј"->�Ҧ�m��)l���,���?7#b����]��'�h}�~���{AqmNB�x�_bҤ*O��?�Lp����NV�}_�{�(����r��dȜ��џU$�gvg�nڏq�Ѿ�퓲���xji��u���	qYA ��3���X�����;��^Q��>� 	:h��Y�Q���Q3��b���Ё��NI�rIx;�EX��g���+�0v��~���}���,�5CL�;���?[ �Ҧ�m9�>��8�A핞�7N�oR����z� FXK\f4[���l��u5��3�T2n�c1�!������įDwE��Y6�"!h��-<q����#9��{�j��Z���$t����!��օճv_*}Y����'M��X�L��WS�����
kB�A1�7H����9:6�bW�<�o"h��CN6_�y�=ZH�k"��vG��R��v8�]W\;z�Z�U��ǩ��7��&Χ�'J�$��\�\z2Z����6�+���L��G���6��f��C�DY��R�?{��,r
�`K��a,�V��b"�S	?��+�-�+k�� [3ȸ���������,[���u�7rЗ�8|V�����{���r�o����W��Y͜���X2�����%�uG&i)ԙ���B���R	>�|��4e�T]�B4w�q 9��lX
KL��G���
_���e�r�8'tU�Hye�o�ZDWz��h��v ֑x����	��>�i�X�@#��&�J�+K���r���a�<#����J Z��Z��JX�k�*�}�&������dnr`��;K�52���ƺ):���˛|��.LuJ��u�Uz#�M��=�cڹR���L�Tx-�O�~���|#; KA�"?��
��^L���3��L�f`�]dy�L{�M
6��v$��H`��BE�f������H.T��L��ݚ��c�奨Xp����.1ќ-�l#�	DX[�_�w%�K��"��|s20�~I�(m��v���������h�����^!#2�*Y�V� #�3���H������c<~���	��Ġep�)/DKRr����Y
k �=+J�J�t���[�h.wH{������	ͮ�e!����-�U�L��Ż�ݞ kP�eޚ��fYe��.�"���O��XFv�����L7�A�lC\����H�����-��O��+Me�� ����rN�g�¤��N�;��$o�˚`�R�Tʎ\��:�����iO�}�w��+Ow\�T^�D8r��֬�9�_�u��Ӵ��p� ����ך�]�Ybs�H��s��U����~���lg,q�ʣeZ�%}��W�1a[+Z�A���Z����)���f��iQ�R˻��v��'*���r,ؤo�5�Z������k;"M��X��e�U0K1�>��|HNĬ�3�^G�3��[�5��1��ŉOP��e�}���7��5~X�lI�3�Y����X��$ʡ��]s��la��`���W�d�0���&"w�Mv�wI��p;a��+��1�����97�s�iu'!�Y ����.ñS��������fQ��	+H(�O:�?�Ӱ���B{���]. 9?�y�!L�l��jK�pɗ%�P@���������6���KU6�s�?���,��9+]qi�]v7��Z6H�|��ǔZEz�S��jI������t�cRrԚ���|Ź�X��܀�h������*d+��Z��ʾ�(F`T���69�j��t\�A�!�E��T�[���'-T��\D�t���-/�&@9�̴`�^��V+���R�� �����Q���ƖP�?��b0��əb��;E����#
��Q9�G�e���O�K!-W�)�6L��%����������|+w�N����Jg�A�R	k}�}�hۃ!1
��b�,����O�sdE-O	Z9��h`�����Y��3b N:t�{����"&��j�78�[9~�_�o]� iG}��#�(�k�Y.^�%6��)��o�����fM��_����'����6����
�7�� ی)���"��K@�CSS3+�`ϕ;y�����k8��~կ�-��ꝊŅX��u&�˃�e�6�~�*`|�B�΋'���,�g���z"�v�X�$�O,�m���
s���pڏM�W7��ar�Aؠ������U�"����p5�bz�.�����"��r%XݮEK��-s��Ӯ�g���C?&�D��V�|!c����b�UP����I���f|h�孵1�����y񋸫�;��fM8��O�5�7Q&<�O��$%�;�z=Q�ez�p
���Q:.� ��:U;+	�Km=)D��9^�Q$����۹�Kr�8�	k�S��t��5�md�&�z��A��;�5�(TҳP$	�`#�6�J�n$�y�R�4|
�j���e$�8p����TQ�淌�?��D4��fw�޽TKV��|&�O�&9n߂eXO����$Uw��Pi_�T(�Ҿx�葖N8�[�}r�,����q����x�y��hA6���dЍ�_ћ�%WXe�'�����5��c��P��f�A�#RAR�L
�&
��#�(8x��Kم�J� 
��tk���(Op/W�11�j�g1���9�y�����Ac`�G���k8Z������ɂ�g
/��F�Y�������X0B6E�*ƣ��l�#�A��N�oY;W�cNn<Q��_m<%s�f7*z�T�3*��b8�SQ�o�A����.+SZJ���$�{�]i"�ͺ� �Xw�C�gF4Y��L�R�B�?��Pз��ի�Q�����"9x�.���;�����Eę�R�;���xM�v���@^�Z%Eg���\@"�scij����A�����]n�\�R˃�HE�,֙�;��Wޞ�sA�t�<�{��t�vh�[`]cu�����0$��w2p���_r"���~�3��@�A�8(��T N��-�7�v�>o��=�ZD�9@����H��?�r�J�p��c��b��Ə����������m�V�@�%:saz/�?��v��,�e����=O��ҾY�E�8�2������:��ވ�1����e;�<�&�]��k�g�j6k��o�Ȼ=Z��[�����ԫ(A1&�6Yv��_~���q��(q	����zl�/m�.b�'C��Ǯs�h��R���h.����+2��ߏ�<N�姈u6;����(Yc����)�dY������X�$��??��� �c%����Y$K�·Q�����0�y�}�y֞����l����+.8�G��حd3̎�aa{Xق�Qk����H��v���&��!�lK�h�7?ή������������ſC�G�܁�2I��H��h�pC 7��+��u�a�6xX��x2�m'Z���WC�O�H�V6�����z��@�)���������<�i ��9t�"c�zO|��-oVE΃v&^�|{�c������f7؜
����?8�տ|�o�
ؽ+c+61��l���{Q��$�l��Z�g�,B Y+=�X�N�a�>�x�TZ#w�2*�@����b�S�o'"V�{>S�������Q�ءZ!�9@w����x�*'�}�aMV}Y���8]6!���ŗ/��X����`�������]%��K�1�T�E 2r+���]Β�a�Є�x�]?�8*Dȥ�cw��
�J���X*�k�� �OE�wr`[�a���FE�Wx�g���5��FX(&Mw�r�&���t�
�?B�4��o8/���e�@�d�|��'���Rf� ����
JT��X�L.#6[���=���=�_�ìv�R���}IX�� 
)G`:0��/+a����\鷈�R���y��D�@Q�81�n�_N�cp�g{,d�Zᩐ�>Q�+	���C�;f��~�-#ώ?xN���} _�˱R�~`��:�7��bFg�v�B��
f��'Cᑦk1�k>�!�v|x�l(�T'���Q�L����N�����*��d�xq��ɿ+����U�1F�\��m~�P�=�ڗ�?��w+ "�ޓ�����R��"�j*K�[@���#�^afgXΛ�Lb��h^ܰf��� r����R�&"_��a����)��JGk�&��d��g��u�I����@�r|nRa�@e Wu",�k�������$O^�ڮ���Û�u�Y&&Y��I@���b;���c�R�h��y��>�~�P��2��v[�Td����ѷ2#�M�*
���P�����UϗY�kʛ�k��8��u�{m�~$g�r��T`g�ѭI.�@��_��'�Iz̼#$�@:�5J���/)i�Q�e�.�司{�s��<:��XN�� -�߬����$o���M����mN����~S���'�&H�{$����pG���x.a�DI�F SbN��{uy�C#�Ng��dJ����3ɂ^�.JݰEv,,�b�<}NTjֿ[a_`�%,���&�3�:�����*�Y���@�_�i�ݺ�&sN#�1"����kq����H�&�mA��Z;�vU?���}�>(K�ڻ,M6i�����iKߐw��e�,`��i�|���1�F051} 7�g z�?O{E�����M��]������r���͘ҹ�~�9�H(l��2q��8��|��������@�t�g"S�dm���Gз�r�w�z�X��*�q�v�/�#��%Ȼ���L�Q�v�>֧������ t��c,.�gA�}Ȏx�ލ�uJ�{�W��U��a��/��W���$td:?��#��:e��1f�r��ؑ#�u[�GK����v�*�d�Ĕ)I�B�>W|p�/2:.W�{�u��2��8�H���v���:��-H��B��������I����x�(!�
:LA��z�>��<�e���&�s��������� �l�a�'nM�ܬj�W�5�	�	@B�Bz~��;��C#�8�J��YD[�*�W$���������0\�ή�m�#
Qd'���P��t�[K��_)�N�%�1��O�PZ��� HsEQ�#��'|ҳ�t�����u�@����t�[[�F�M��;�(�:y����Ԃh�S��KS��������Lj��[s�+/ ��"����5"� �n��\4�?_���hԑ��2�+�WMW��wW��;�yk�aRz�y�%W�t}�F�n4?�PT'�a��k�*�E����j�'�O�I�!1��@�xeQ~�Y���&FR�P�ϓ�cC���]�')������������!�5���c�5\���y(�k{��;$�NCl��u����#�Жp��dA��0>m���#�ۿ�D(����R�	l�bIZ�Y�?��h��l�מ��N�F�S�w�!P��sgλ���I�������
z��P����������B���[��$�*��RfOo�$vO4s�d�{��[�L���}R>�X�����{!��k�{�#��4�Y���Y���/���eVs�"��⣧�P�u�bs[��͇��j��Gn���#��DC��y���!�y�aH����hJ�L�r�h�1u��,r8K�UD���!�)�w��X����l��B>��1�u+A��D����N�$���Φ�3���bSt�x�p)�z:G�;7_�䋫�i�}�J��=�WV��ڣa��5!�Q�7R�Y���JX���S���Vux��-B�n�L)�.?'lՐ����XQo��ЩRߙ��p�/`���3܂)lPp��	4����q�S��L�
�/�T���O�.��P��Gʂ���
(�]�ϹO_*f����F)���Johԯ����xb��n!w`A�N�R�XlX��F|��5u��:X@��E*���0E�U�$�T[��>o�ԝC�	���_�� fN��r:=�ƎrWГ�(*:�V�~�ϱ�Z�T5�T�
��~q&I���ؿ�a�M�ޚ	 �(�������?�+k�B��<���jG9z���]�'4�:�e�$�ⶱ+FwT������$�-d*#��D�X�R)!��C��rC��I/h ��;*�f�ۨἙ@��Zfr-˶zFH�H������S�P�4�}�xc��[@��:fg�zU�-�爏��P�&}崼3N]���y&ҭӷ�i�?F],_0��Q]�o�؍�/5x!b�u���S�ς���׎fOE$.�?��~�]�ӑ�߯[/�S>-I |l�����_j���pͲ� ��4���#�T��3.�9�9_��@�/�i��{x2:�5���p���c z���Ѕ�l{^7,4���z�v��J�in*y�A�ǈl��d����֕�}i���㍆ϐU�
*{��z��`iK9
�m�o�Z�ą�fs�W����E��������x����S
�yһSV[)S:�M� =$����<���L���Z�r���dg��b(�U����ڞ��٭ܝ_yo+��b|(�ܛ�QUfu�������JN�`�gqFm���Jzv�7��n}���K-4X�Z��6c>0+64���Ҍ~Y!��s�tb�	�L���#�y7�(wD�y�8���sYLy��+�J+r�.2io�
��-\n�h�i����T����M���*��+Q�Að�WP�V��&�si؋6�3�AbrTRbFlGE˫�-�s*<�z�)g;L��Mv\؛�ARP"�	�{�,?��v�>�ɶ
g����y�;$G9�r�����D�'\��ә�Uz��L!����r?Z��;,Cs�.�q�Q���ۊs���
?~���A�}]�F�y\)����L�٭�����B@?�^����w�t$L�Iu#�����������0�������
Je���8�8��$�N`���D��Ū�å��K.�w/�T{��K/�S��&^�\_��圿:M�8��ԩ
.�j5c<���7��,���ދs�ro��7��3<���]�' ������dCb�&}�R�۩`�?�HKP��x�A*"��HS��Ty_��o��8xw1/�p9��M&}\Lj����{
�m�Q�l��,��A�C�\��ᗈ/�Q��	��<������T���e�Y���6N�d`<��u˼�i�~�����b�l��2l8�����PTb���քxk0���LSsarS���Y|Bk�W�a>��F�|w��� 1���qS������߭ZG��G�F-U0�V��Ń�l���ùX��K�Ҵ��Eq%V:���jߧ����+>�@���{���IϤ;N�_��G?��x��ԟm�NJf��I<�� 5˯�e�~���������>�;�?��I�q�����H�"J_�Ł��vގ��ſ~�r���X"����w�0������ºe^�A9Uݲ�a�w9�Q�K�br~jD�~�Q����v\��d�˪���t�F}��+�c��\�|)�Ŷ���f����|�����Q8�TO"���I|�p�<��G����H�E
:&���&��?�^U8�O�z^�9>�>M��Nv�u�e�=K��(SH���5d�p:6_�v i�O^���X,A�baIj�b�g�?���ө�<'t��L�H/K��(��' :E����7v%�+��ܘunPYr�~6kq�ᢿIݷb��{vj�>�6���Xllw�A��� �m쎠��GM_'��?�_?���{]g_������+	�u���0����	$�zSiA�	��X�`�sYX+�ǯs�Ϥ~ w��a^��<�I�%�p��7��Yi#MS��$k��ޗ��5���?�����n;a2�111qc���#9s(���;;��%f]jW ���ܥ����e�|����>�f��]�S�Į���N8>*�����y��4��>2�I3�Q~O)P+.�P����%
�E?����ӵ�"� ߗ�,��g~N�uq,D�?'�m�Tnl3Y5G'��o].�j����w�b.G�fҖ�����çm@���P������ӡ��{N@��[eMM�Bڎ^�,��3����]���·e*|�s^#e^�m(e����"���"]T_wz�4[�L�܁���߈+D�<#���x�H9�4��:���$|����ݳ�Ҹ�<��o3O��K�E�ۍ1[f��g��Z�&oTnϸ<�T��cU���N�W�x���J���8V
'בQb<nV7c��lfKLm��{Ă��F��V���'�͞��W�O�oI�Rԓn�$��5���ӞFY�>��	��y2��d5c����b=��s�]E��e���������byY屮a�4���6P��%ft =�){b *�_��:{�⭣]����U�C^�͇��$=r�Ҋ�8ïKvCr���{�c�>oɔX���n�U]�ý;+�m@J�5k,D�N>uylJM�O�칹a��,omÑm�����Ny��J��K����y���`�`�.�埽\D�+t1��A�Et���rp%?��l��Eb��/�n���tT2�-���`5�^A��S)'��V�"�)�;�h,�İ/��6N �7.�,!��,n���GF�)�&��>��W��t����';�A~�}��o�Q�ƽ��3����D0�W.�ADBr� Q��r��aQßƳA�J_���`D�Bۙ��ჲ ?ηo��%�3'�?	%%G9��q���=�Hăf�#Tߺ068b�[I��n�#��	�\�D'.�9X$��cݸG�p�����(:vsʞ���y!�*m,:���z�=�A�V�f�FR(i�q��o�t�6������,����PU�֗�ϐ@A<~~�S=&`9?��_���^Qn"p���h-RD͑A�����Y��c�4�kק���oA��;��E��f|q�0�i�!���6����?�h�I�Kе����[���6��X�6���%g�r�Pv��j�^B���C����@�R��B[+N����3�n��J� �:�%��ӭ���oor������B�c�Rs���0N�V*� k��^�za��v����D�t�>��	�9N�,`���K� �&�$���5G��hH�#���'K��2�����@��3+P�p���y�e����(v,��o�_���¾���r+��/��X1W�#j��j�>��k�-Q��)��1�N�y�aA_���:�m�>���׭(b�B�E�ܰs�9����W���n�=���n�V�lg��!��yeq0�����hrZs���_b��ba-�guJ�wF�Pq��W�r`Ǫ�FB�(��������<��g���� ���dU$����c������u��;��u��JR��M�w�fCA�]�2�B:hӼ��V���g�N��2C!�S6��R��rz�݇�6/��L��s^�
T:�t��q�TC�/����4�8�ɷ�#	�{ycY�L�ܴʵ���B�o%=�x����y�a�_�gVz�	{��Jq�&��76%Au��Γe�f��*y��+J����ޛ�C�v��/�R��"k�v$!�v�J��mT��'�蝢��(E��}�d�:�Pc�f�f,�;�K����������������s�s��s�s��^���_���J�����I��ƴ�:z�U����7�����q���!m0D��ݮ�蒖��c�m+����-��7+��1�+u[/R"���7?J��9����������r�L7YU���iV3��(9
{���eK4	ӑ;�j[�@���gÖ��}����Ӛ�E�]j����Ұ���<�-<��w�p'�$���	���cac#c���x)ϣv5+�O]jf�X4N;0�8���29�۲���ڰᤥ�y�,%�S7<��M�xX6��s�1ګ|������I��שּ������W�����ː�&��r�]#^FIjGc���s
����uι��׿�Ե���Xf�����s�d4wE��g����U���1�����~�~�yc�9�W���skKNn���2c�pu%�c1�N�HA��s?o��c��3�*�m�z�ޕd�3�,��#�n���>��[��[��b8?z��3�ĉ\w������_l�.f<O�g���B�/|���M��۩���췍������ٺD�ܗ!	�{j� �ӫ6�Q�NML�9�_�Wr�*�f�is�I�����]��D�U[qf2h7��c�"���@��J:>yCx�`����9�/����.�w��pS`�>�G����`b�C'6�W���;�^�E�Z-VY̭�w��JF	=���9��\�`�]���'��5έZ�~A�����_�T�|��o���˿�[9��f��+�T.�M�y�^���%�mj:�����cOC=*�<4hǚ3���b�K������������ ��g�W?�ѬΝZZ��(�)����"�o�-K�W_G���b�鷞�O-�>%��n_O.��y��.�ѝ5}=+u�y^�/s;�d���˸ysv�Ȝ�7G�G�W���S/�d
b�����oR|��Zj�m��9���+��:|�Q:-7����_H�-lq��~]�ċ�W�_y$e�L�ڜ�Q\�Fx�=J}z�zۅ��� c��Su'
5����7_�q/������>/�� �
�L~�O��V|/��I�umEՎq�1Z���|;kM/Znuk_ؘ��R���Tt��|���<a/LF=g�����0ۻw^�1��>���mҾMR;�ʙ���q�C��Y�22�a�̤ꋓ2����Եl�]U�X���=Mʜ�EnSq-%�Ѷ���%�_�yP��~p�h-�zF���
�Lb��N��	|�n��^�l×xb_�I��;���خGR��_;��m�2կ�%,f�i���{����ޭ��n�������օ6��cY��2L&J��!�}���i<8T�M�΋<ZDiu�$�Jo�k�)`�._����ܥ;l�n�OK[��)�O7��X�g�����D�c%
��Ԕ�{
Wg���UZ�՞�zc���W#{�9�ch�������?��s��L�֙z����C�����<�ff��u~������|�$Ffc �hڴ/�u����P�z�&֟�m(���)��9ɛ�ǧ�Ǉ�J7*S�+ޅ݋�h�­��g���Ͻ�e{�BOY:^�%�D�4Pƽ��N��}�1_��r޴�X����E���*�u�D���&_,�w%s2F�G�:�:�ޏ�V�H�+髟�[5��>|e���dw�Aj��)�8�[�|�O����~�����,+~�7Q$���/0�
Ͷvb0Z�F��cV�ݯ������ӭ�~��Ԉ?�on��B}��i�d\�r�s�q�}�E%�i����4��Gj����W]���[Bw�����b����D8�a!��5�v��w�V�#��hˀ���}:.Ǘ���Ɔ^U���4�J�}˽�.��)�y\�@�\����p�(F�1ổό�ֿ�e>V>0����4��묤�y��d������O�υ�=
�>q���zR�5��nP��zV��۝h7���S	�}�KD�)�ǧN��#.\4DT������;�m���|[�@�O��f�ǋ
�{S������?�A��xr�u�I���~��Ĩ8�����p�۾�z��и�b�X��l-|�}T�Jyf�\�(��[�"v�R�vD>�~I�H���x�k�<�$�PT�kB{\M���B�]�N{�9]5oiRR���YY?�a>^#���QL^�N�'M[�E]���:�:�g�����6^oZ�r�y�'b��aY��s�.�X4�,}���ihbK��w��y+��n|�>ʵe#�ofO���&�a��ΰ{��>h �L�>�>	E�w���n�9���6{�
�o�3�x�L.��wv����7GDb�]�z�a��n�h��3-���΄x���.�/�ʳ��jVa[X�.�<�,&�q�	����M�s�{���s�aq��a���}Q�O*6	��n`���T�d��5 ���WeW�
�	�<��{�����ۻ���g��Q�y��p�������[��[��7�3�G�_��Q�*��;�P��_���z�s��g�C��E)Z�Q�o8�J��eS~�Z1��o�Ck��n�NML�ۅ��v��]�d�_y;��6�SnI�A��7J��K�Cj��1��sԖ�|.��Yb�y5�"߃��__�ל������O��Ӊ�R�#�E��Ϋ�ʧ�������i�ī��e܎7�b��Mc�h�����myg�6�7��hR�D�,l�^�����S�l"��j�_�ϳ+����&xwj�g�v����ô?am(�`��	�]�񦀐�}������ߺ݇
]�M�����ɠ�h���g��O�8��+�?s�z�ݪ��9�ߪE\��w)��9c�7�0��ϟP	�O_�i��ƣK$o'^xh�S���P�zN֮�|o��.̒ߥxw��y�\�%d�i�H��/و��G����g�6?6�b�.SYO'����wj����+r���=�<�홱�K�-�Q�O���s8Ɍ����Q�cKʳ`�Nx$�g����������U��#c6�������ʡ[����v�K{L��)��Mt=���܆����$���ك0Ҫ�����j�ɟ\�;+s�b�SG/
�,��mU���V`Wf�������>_�x���iv�.���_{�V��Hm�K>����j�qS�����+冋�4t��t+�Ժed:�w��hy!g�'l��JÎ��.v|���wb�/N��11�q֊����=�Q�6��o�vM������ҷ{������&q��^q�iDA�8a^��>�������և�*W���I�T��k袘��Ч�,l������Rڷ9����i�&����wO�ND}r�{>g�9z�i���b��D|Xe��J�7�=:��/jlx��!y�x���r���=�7�YR����/(�������������\��ϧ'�vPW�����=ee�t�x����i�~�-&��&��(��/�p������ZZ���9���a؋�k�Ԣ��͙뿽��4/��h,��\������'���VR�Q{/��Z�IJ��Ms��;.��^�)ǋ�>���c����g��]5�ʯ��L�c�U�>�j��iv<P)��_;QW�n�?�պ��n���%G�I׾���r�iK i�����}/VR���C%�:s/����x��1g	������ôiK�h�/�����oJ����)�X�9:u�{u-v��pF�s�{Ea�7Ocٚ�9>��M������]y�8a0��#L�hʱ�o����NOQ'o��.�����S�z&P�~�2]���l}��F>��,��:��S�W�7�U���u�V�@{!l������_6C�+z��<�V�UⰧVR���h��ܫJ�B��ˏ4�q���|0�m�aȾ�ݦY�Ǆ��)��~sNȸk�(s�Yu���+���z,�]���|8m5K{�H��Z+j<C��9���n���{<M�X��>���Ǭ�W?)in��]���&�w�'G�e��äx���;�rb���!;�,�{=l����}�@�\�IW7�}��㇬�����F�����SҿL?�n�5uַG���uu]mZb��.M�9��T�zj�f'9�^4����B���P�/��x�����I���n�@ �Ǒ N�2�3iM�]}��l�UM�*q�Bڇ��ENF�:�{��o[�-m�j�j�~D��l�fzJ ��鋧~�+Z"���wv����w��j�7�#� :�~�a�Ah��i����D�+n^��Cw�Y֩�����u���xmh��[�D�o_�ft��H����J��P�X�D���!�~;����Ry��{����M���ڔ����'��G<�Y%�?nlZsm�Z�'�\�j���{�Тڏg��Ҏ���W�?nM��ˇ���yn��6U�vEF�B����^���T��?*�>ǣ�&Ls��D��ģ��'��`j2���g�j-N��u�z�\^l��+�0Jk�����n���k&���7����T>/����k�e�m,k��*�a\�^�w�~��yo�%�Fn�K��{��e�<N�%��O�V4��n?�\e�d����P�=��6i�>��,ǔ���#���~>��{�ޕS�#�G�G�)sJiM�m�վ�����ΩՁ�Z7�Y]i|?��v���}oXaY�9y��O���u�7�m%"9�G�����<��ϧ�N+��t�MN,ʌ������_��#n<��l��N1�l�ٱ=p��*OK.�8I�y�$U#��N�<�ױf�i��*��oy\�5M�s	�~<]�){\�t�S�C5�uO�U����㭀���C�yJ���������A�+�ۄ��=,�_�r8e�v����q��Z��o�y��V���r$wqװ�j�q�'��,�\T�I��\X�l�|Fv���ւ�L��.���z�Zb�r�Q
ơ�g�m��nX���9�r����m�����+�]
U�t��xS!�v���y�g5/*��ٟI��yɹ�|܇zi,+�'V��q�}�e�Pv��f,����,��`�Sj�m����;>7�~c���MYⷹM��~�(��z�������s����S��j{P`e�ʛ��)G���0��=\I����"~3�n<b݌�3�L�tL�*	��T��������z��\]W�<�(�����^�������?�:���xH�P�u�T�V�*�oK6��T`#u���̭�:�m���h�]9�X�aE:/q��F�grL-��4яK����'X~�����䕯�+$j�~�<PV`S�z�巀߀�E��N�\�a�g{&I�_�ϻWǗxui�L��g��Jq0S����l�!*+<9D�UK#�B:pz�����}�v�ҿ�<�:�3�c����"��e��p������_Yx���XK߮�����g��iK�?����Z1<��[uQz����Α�ŏ�kK��iO/W���ݷhI��v��gf+7�T�d@��	�~��4oQp�e����E�n��Gm�U�X��Y������d=m���✞�V"�QV���νg]@X���Uz��Zr�)[��)�ȁ�h�f�C��.-�m߼8Y�k΃K_%�ww�"�'�~�p�d��C"�b��зCw����*��/b���w�Y6�����V�S�g�X�0�حԾ�*w�����W��H<U�#��wa�;C�`����s9�F_C��za�����n�O�}�p�V.�Ӕ(�T�YwC�?1�E��oV���9��+Q��48LZ0q�	��֓�U���#�G]w����*�׾G&X"���󔉏Q�0h�Y��S8�A:����TT�ٷ��<x���C�o�o=�}��C5�SQ��9P��=	��*_�<;r���˸�����j�+àw>��+�vh�?V��Sn�>���<�\0��9����u��EI��}=^�=�cѣ��︝y�?٢|��`���w%lҤ��N�����,�A
۵$n�݌��94�-qx�S5�p�BՂ�\��&���W�`�Ȗ�m\���zk�M��O����}�D���o���Q\wZ#�];'��8��p������V0�z��{U�Ò���
F<Vڻ��m�݋_*'2߯#�1WB	�%_䵙��׾DX��>vŻ%w����q.�J�Ej<6@��y㺮*˛~���^�#�x��-凛�{�3Ft�ɒ]�^.�崙V�e�IR:Ń�Ld�:<�j�ߦ��r�U7�!�պ�J�asS�q��7��?�xb���Dq������o?����݂�'ory��܊�6r�I�%k4ɍ�D�x�MA~��������_a��d���ݝ9��5�򫬞��c�����t��^�Ԏy۵�ڪ�:���H�Մzm����5]r�C�X����|]X����;<��>+������ɟ�*����Z��Y@kJP?2x����Y��2�����,J:�� �:��?�t`*-��Ӕl]�azG�`[��K�&M���t��X����O��͡��ބ��=J��_rM���FUKb�N-���?�T�`?YW���)p1Xb�?c�ܟ3,���g������W�NW�j�M��'�.^f*(�w^�?���XU���k~�)�o-�ǎ��1,O��1�ʛ"�b���c2�Q:[r�{�h��_�"+�}Mјؘq&Mc��-�a�kQ��N�[���bsE*��o'������|֦�=Uje��S��8�����his����֕�W*J�
�jj�z�~��d�%t�6���EG7`�<���&�.��bYLx2g�{ұ]�:��/������7)P~25�Y��u�����I�������;�gH�z4���"~�s���?�jv>��#��G���n4m�xt��������\�+ϥ�9O�~�kH��>��ٴ���O�5��怟Ϲ�Jκ�C��E�(o��mO�p�b����V�<q����?�����F�%��.�U{6�-j��{�r�M��VEo��{���-k�)ɿ<����[>s��T����x}x��B�BE��&����oW����\-���l�C�j�{�0�],{Q�&���%\�Z	�d�Hϕ6�n'�難�MJ��!R�/ރj\ZgI���.�s����s�m#+�O��7~�i9��c���h�/�d�E�CԆ�^D���N��i�ɋ��8�~��7����\W���7�\��b<�Xy��
N�v����מ3�A�u>�Z�ɣ
�����)0��,=h/ꜻ㜤�ܛ��~��-���:H�a���1�[L9��;����pFzK�c�=���J~S'��q��b\�M>Ƿi_i��&��^���R��� �*��yi��F��Ãu��i#6�Y�����l�=�frTQ��;�\�!x�/`��'�؉;?�o����F2��W�f���d}߅�;���&u�|J��RL��'�|���N�k�kT�H��5V�B��o���{b���k�+� ]Wqo._q�<�ڻ��Zb�O^72��S�-B�^h��3aRV�|u����ʊAOxP��S�4y��b�L�"�l����e��#�w�f�O��xq����hJ���I��}�o���]�� 	�D?���s�;�OZ<L�~�W����+�A�ІҪ���v\[���=��4�Kw�i\>Ns�o��yi�k.@ӺO��0�F��=�t�E���Bs��q��OMmi:Z/�ۥ��g��k��S�_L4�|�L^��k<�"��r0�͡����$�P����H�.��&����x����J��-YS�}�m�5.U�K�	Y2�D���K���/�W<�������o��
��{gB|�$I<�?Ё�S�3��[����Q�ɱ<����]�k!�1s�c׮)�u��x|&���&�u�V��s3�&6��L�5�q���#�f�ՉG;"�]�w�T���M�q٘�>�w�H��k���]wr����CVO�>~>����.��K{�2��X�����N�>��n{Ɔ����r�Ǹ{z�a�4:���*	���)��&��&��Ð������h���Ӌ����R����oL��?����1-WC��rW`�O�Fs-��7׾�<�H����r���8�|N6��vO[ p
(䍄�K�pD�*��;�n���\������3�vefO��n*�����蚉$�49v�t�d�c���Ѻ����[��������<xpN7�X�/V���[(C#T��ڏ�n���L��е��Ѱ�\!�R�B瘽v�l�&�����w�Z1���Jo����菻����%��_�'E��S��	����[��(�*�V��5g�IP���y��&/��W��)�n;���e�o����m�"5_$T_K�?�k��wd�½w�^��;v�����.<Z��Y����M�+��l&q��K?a{7�kR��:����Y��1�I�B��W�_�헒W����Lm;3�>f��n���wK}���KJl���Y���)[��OM���s�2����ύ9%p�����s1�s�0+WVVn��e#V��8�K�Ju�Q�}뽂�jw.[,��>�l�΋!�:&����ȏ��fq�CAwf5?�$��شcC�≟��޶`o'�:��6�����P��/���h,&�Z �5��K�h���xʌ�]�񂥼��o��<{*���JF�A���鈸3R��0���0F9��fDzi����T��1mo�,E�*�B����b�^Y�n��D����{�`�8��'��cq�R�)9!�ܴ��/���T,�����Qj����q�z��1J:���ȋ�M��Kz�J��MZF�b����J-5�?�M�3#E�1��<������SW���ˬ��W�Ͻ:\5�9�����k�W�t���f���kxTv}Kh
���1��������1�|sB�U��I	�ʋ[�4e��܍����ȍ������,��ӵ�J����X��0 �Pvq��阃���ƈ["zx���s��n�\�y�']u���P��I�q��;����L�(����ٙNK�C;צ�S���\*�x��ZX�����R����������$N�+���M9�k=���x�'�w3Ft
���Y�Z�ex���:�E��F3o7Dϵ�0�Aܥ�����I�z��_?��1ʞ����.�+��.⣅.�)�N�n+#.n�k�,�@㾯�όj��PFTdh��0������e���u�bo�3ք���u�1b�GtX�i��e!ACؠkP��H8k���� 
y}xb]����`���,��fj4���=u ~�#
�O���X^�P�d�F�.8_�{u�Y�������~��t��"�#SA��IvF����X�kӛ�����v�e���<�j�ؖ�(���1�4?�����Ώ}L�"�-��M�<�zW@67'n�}c»����)=��*iکup�x�:')�)�I��3Η�J�	���a���%*-#�5|u����K���
�,�.�Fë���;�0킮o5n�c������|d���=˓t�!��?��|4=��d5T�n�ƺ��V���5oL�FFds��fh,t�Do�_`�;Kk~�2zk��,�s���H���&o���u�Ē���Z��0'4|^�)H#%-܊wBesٳgy; � CA{���i�&�[�b��@�'��s���כ��|��=���ҏ�<e� V�ЧI���;���ٟ���t�3��$��J����l��n��j�0+��^ʈQ�>�2t+��$�J�#��CW��s_�� ��D!_����=J��Ҁܺ�+4�Fޙ��@�J0$ѫI_�)8�X[#���Ǩ��}1 }��d�p#�h�ff��s�}��I�*$��e�c�SO%7m�����l01N2A������涊m�sb�aa�D$����ey�?�4yH���N���?{�0�rDo��I0�m�vo�Լ�*���(���g��Q�#��W���܇�z�]�4��M��
�@|]��1�O�����ِ�جB�;0��L����HK�8k4�a6dh�� ��Ak�� |������ȳF�T�'�����Sv�����ќ�h*��]��Dl�m X��/	����k�1�ȁ�Fx���#�ťqi��q8C�hߧƤ\��^}*|q��D!#�?߇r�ء�ɇ�Ih5�۫��uS���т�U����az�BQ5T��S�6��o&!���?��x���>�9彣�Y]@>:��1iD*��Ԇ*;B� ^��E@o����s��t@+���=Ϫy�c�V�mձ
�a�ֆ���lH&nw�sr"GtΜ�����0�fD�q���X��vd@AJ�s���Bt��S�mD��[��*}O����e^����~d�� ��@|"bEY)��Wֻ����YnS*����|`1e���|r��z�6R���lj�W���8�Z��~���������X�s�<�{��:�p'����Ǆ|9�5�8�(�R��hG��?�^>�n�K@��{���G��� ~�T��+��)`�"Gr.�aj{�Ėd�i?}YiF4��:�}�ⶣ��!�[�f�}o�P(j�[oޜl��P(�P�3z�=�`ɢ	r2�]3��s�#Q1����\wv'JR��l{� f�Y	���b��/��O���wļ��j-�߳�l���٪3�@h�V��!�#橭V�>�Ě�}����=��6�Iy��ȉLZT�b�w�	A�ڣ��Î�x�IpP{,.�(����v&�=|8�-����X��J5=�퉡��6�n>�����5�ak��ຄFF��ng�=�����Mǭ�'��O%��)`��ec��|V��#�'I�b/�x��񷿞�'���D�"L��{{�'����lD�3����S�<vsߍ*�j��ԓu���(��ܩz��+U�C�?��P����폸u��G�޳]�JBv��H=8.����}�����S�A��9l>�D�<�w\-�t�#K���������"#��S\G��Z���=�u�d�r~lpI�����G�aO{��ͽ O���B	c���@��o�a�d�#��j��3f����}tƿ>vcVaVaVaVaVaVaVaVaVaVaVaVaVaVaVaV��z�?
����/V��V�.ۯ"1�A���^�;, ��w��k���:�ή���:�ή���:�ή���:�ή���:�ή�+Zw6D��(��t�|��~�vv�]g��uv�]g��uv�]�/\n���׻ �_�2�ή���:�ή���:�ή��6g^����\P�g�gbE�3驖I�Yh�&��-iJ�W�������*�MƼFtc�=v?�u��k����_���j}�bh����z�Mm|����l�g��+��mg��50k`����Y�f��50k`����Y��_P&ߘ��d���7���|K�<��-���(/'��v7���2:������wb�wI���|/����r�yc�
s0ڈ����	O�w:�������ʊɦ|^orDor���?���B���RxE|�]�,9�:1y���C�)F��0�ɸ��?��/��,��9o�FM��:i����i���~T��b�\#�{OﱱŒ%�e��'*����0�'>\ՈY)G=��-�H�X���I�*�������3T�W�| _��WQ�ĤFA��x�~�DRY����NL����jIc�b�Z؇�T���Pu�z�&����X��HN�b��е̠"dF�,*��r	>�� T�w���pib9��nvb��ɸ�_Ȱ2�����&����߅?oUC�,E�0����y��|�퉊
�󏼃%��Ɵ>��iQ�rE_��(h�ہ}����)�7���|P�F���`&Lp�rl6t�P;'I(���=�`�E%��~�O�����{)�X�](_�F��f���N�r��\��kޝ;1y'׼���2J�؜��ڠF�ܪ���&�a�np1�/ӡ�1"�
�n���'�Q��Ȱ�,M��l���Tx�(�����%��>���?�SL�u�eQ=g,�∽���qΑ��Q.��!���TB����.��$����'S��R@ċ�	�G�$� e�B��(���Xi��sl��w�nF HB��y3ԑY6�}9��t�O����g��%N�* Ჷ�s��n��#��+�3�#_~���>�3 F�#n�Cʼ��<�����]�[�!�`�𶙡0����%`�O�y�ϟ�d(#�5�9|r�)�3S�?��Kt�Iq���nHQ�*��ݽ	�������8TN37�D�!t�7����l���q��p��~Ri�yG9��Cԝ�I��2'�*(�Q������F�, "r��Vt^)�/���-�����QVe�ڂ���D��%ePbMr�T�2�&
/���$�d�Ex5�����L5z�ո�����Y���Ah���f(��iAI�1�t��oj�ā����/�d��#da�'Ya9C���`)�K'�Ā�5�#�QR�/��30
���L��ڸ��tP ��Ӝ�IBT(��)(���q��t\���ÖL�I����� D?�J5�K'�.�U>1�d��Qo\�+(�DdREPܷ�<Ce��U����� e�T�V� �ԮAҍ֙��.�+C�T���Du�#���w��2��əR�t�֔���݊	zc"lT�:�����b2Ȭ�����>��C��6�s��U �Np3�u�L���Qg')�ŏs����nO�Q ,�`41�H�5� "�5�Te�L���	FʕO'&?ч�>�\+} ���F�L-��"����F�́�-�ٱA�]��WPg�D�VC������98�﬎�B�Q����3G�w�,)Q;<4�ϟ��������IK�0lx�>s�l���������N��V&��57���!��&(7��L��upX�ߐ��d����q� ��>SC�zh��w�ߊ�0�3�^�A㜭35i��12��*]?�,7�����wa�S� q�Iy�3A�v^E�P�2m�;ᝉ3ѐ�
L��͠�z�D1p�DA_Tğ�NVf�Pј��)���qj?�r+���(Cqa?�\�.=�u�M8Ȕ����	���<�F?�PCE��qxp�L+�Mx���H�S*d$�q��������d�<.�a������o\
�#�`ɝ���qѡt����X3tdt�#�6@GF�؄7�#>�
N��J��������ѱ	�0i�DV��Б�R�<�����	�+�^�A;�� :��������ꭔ�V���̡k��Z�2����׆f�<8�C�����:�Q��@����q���KG�A�Aߔ=�L�+��S
�����F��[��鈎�@��}))�a������l�����«7�5���u�'�53t����Eo��a��T*}�����I�����|Vv;x�`�8������h�S�+g~P��4t�I-U��wH#g��ۣTj];Q��\D�}x9�H0��; mF[d���[r��	� �g� �� �_��'����n��4���.�1���H#_[Qa�1��G�Ժ���]zR!�E���O��U����Ol�~�K%B� �Q�����2�5h��-e	[�bOQ�����|�O��>�Z�'BI)·r8n�ՙe��4�_6T��Q���&�9�}����� ��^8&o�N3�������'P����g\���`hC%�}��%P�i3���@Q�l�5�m@ABܘ�����م�l�ɏT��Yd�@����cXLPv�#��CVW�2����d�eP��N�����f��pP�gtȍ�ƕ�����������"��YܸG?��ɹ��?C�S!��wg����J�C��-�h�5�!��yS*���U���ȡ�D����C>�T&���^- �&�V�7���'Ɠ����H	���ߐ�^�E>5¬5�v|�BD	Qb$n������/�|�Ռ��F�r�u'����\���F�y���7/����F�\�An�z����qo|*���$���+�9���������36;�ȫ���p�re_���:~R��D_������v�Ers*g�s����G�f��L�N�HS�D���wKQ�%�@���Ar`���ޕ��Gy�����r.�.B%��3ݐ��?�a?@�o�HmӝI%�t��oVָG��S��:@u���%�� �����$�c&MG����Q������g�~�x��b��"u����
 �9�34�T�r	�����3I߹&��1��b{��w�@��T�u�f��c��ȑ WVQ��19�}���)���:�|~/��;�zO,p�#����b$��޻�=`���zo�z������`��*��,���\4�^9�Q�G��Y�ȋ��1ȡ7�c�ģ�NTQ��,�s'�5h�(TU/�@(��J�	0灛{�I'~��M0|&+y�����>�N���O� ��0��Kj~W��$a�'�L�K;QY.���Uǰt�O �*��~ �W���Z��_3�F��@�x� Jsа8���%�Tu A�Y���p�ͽ�d�!���2Q6�}��d!��O�42@X"��M턽J ��d���s_S�׊��A(�(.�*�^&C6CR,�2l	#MG(]�@2_$�F�ޢA�Yr�0���.i� 4<��R�W�$�E�!+]ڎD_A�;�u��Y��h;��N2��:��]����J��!K����-c���"�!��%%�ˬ�;�ډ�o�{õG3$;2(�U�b?��$F�#�E*]r��fGجQ������߲�BBpݡ�f�:K�&� slD}3W�N�z+~�D~H����K��sI	��^���.)��ώNm�{��=��܈z����F!�A+�Cw*���fT^�p�3�	z%~|�	y���M�#ݸ�tIl+��c�� s����(�q����-�� �����qX'p�n�鉁��>�I؋d�H���2�e3���Jګ{=X-�[zs��Q���Y{AF�A�*�1��L؋���n{�,��{�\��ڤR/s=�HF2M$�YiSK6��#���{7�#{����"�˼{Af����D����Z���)G�"^����\�'��?��"������b��(�%��rȗA	!�B���U��2�f������-FSR3�w��@0#u&��9��߼�$6z��KfX
��RtĎu�&"�:��f�����tC��9�̇�v�._���X	-Qף;@�r'w�є�:Rż�Ԥ��"�	|9V(ƕ�(@��^��IG�a����8���蠨��h�$�1m!����=�����A,�B"D��Y,�l��� �1��/!�_���5��)���|��Y(ʖ����I�e������)�/q���;m���QO2�iY^�EV���r醌�`�����dt�T4���yg?�_��9�~��~k۝Qhs�P��Y�12Y�2w����b�e�a81;�)R�@syM�q0����G"� t�����5�B�`��cq�d3:j/�ƚj?B>4�e��C(��HbO�RC�E$��˭�' v��-*4,��"�hX�Pǰ�)u!��Fj�j;r��5h��f�Є�(C;Cmr���iY~oL0h�\I�����a=8}M�VDZ��Nk;�p�7�S���BC��Z������s�[�B�nPAִ��Kj�3=/���N��9��(�Ks �	���0I,�-u�Hڔ"��8@j������1@�����~b�0��Ajw�!���?>�f� ;��\N�I��H��U&��&�r���ć�*b�~�Xp���A8P����zp� ^,��	�p»Cd��^��l�����^���_��K��[�����(�}/�H#��؉~œ���!�~^*�sA��S��,h��\W"��,-��q�A}��Wd�w7��a3�ڋ׼$W��ari���� �]�"]��L���D��כX{H)��:N�"�.�T�;,sp
�&�#}j��R�Mkp���a/��Z�S�	8�pk�AMw
HW�2G�i8ő�5@J��"�ӹ�S@*����zrZ��7t�HqeM�c�^й(����C��q-CK�h��ʐ��A�l
~[��&4�cI��V�HQ2��6��؂�]d�w�.�V�܏��7�2ut�?��&n�e0���2�g|�B2%\c�[-#�B�3���yK���c���{�'��)�Ռ>؋dx�wܪ������\�^�7�} z�^3<��2�g~�B2�P�!e& W�h���$;���>f�}z�p=�!B�W`/��ؚa�2�fx�^Hw�M�w��e��^8Z*O�L�5��=��C�$��8��[K�z����G��K���83c_�l,A� �%���6���"��4���1hkt�}�YZ*�*��V�F,��%\Y�}�PH.idN&ƪj��&Q���Z>���A���~[ɕEe���s�K�, �����$�md�Ҙ�AÑ��Mn�NɅ�N�#�c��M��c������O����K"�2n�\ko2�[@�����������<#�!	�w��&A���B��&h�� ������jЂ�W��(m���DH!���@�f��3\�fn�� ��e˸�P'�=^� �N�8IL'�j{�n���B�A(�^�s��'!��pԗx���9u���{F��qV��X�c_���I�J��C,p����]�2��B%�b%Jˉ��:�-�F��������z���<Y繲Rz���	���1(R�~��bh�3zWAoٍ~0\���bYxy�37G@�&�b�߁�*
��r���pG�.�sWֳ�����y?��k�O�E��`?�w���rsą���%�2D�I�X
QO���|�C}���M5s*ʅ˭u0�|-�:�0R���ڶ:!�C}%I�R��\��-�6�ؑ^�+��g�Ok3K���:�D�#�B3��Ϲw�Y���y� �t���[��[qcB$��>f��������^�'ޮOQ_��<Q�80�E�o��Zd�+�<�́1�Hx®#�����a	0�+��a>ai-��E�p���a^�e��~^�m��0{ �2R���f��L�$���90!�Wq�4�V�K*��i�8�S���B�r��0�?�������p��'s:��ӾB�T%吡VѨ�-Λ�SH���:$��>�"�
�>������,�H"p�2��V�3��(R�/�G,����A2�~�xH�w����J�*��'���~��$����%��`j�^����
IR��]���� Yx�O`8d0�,��Ӛ���u��Fh8����\�k���[���Dϣ��W����-�㋨[�}�+Ε=_���D&Ae�!��	�P<!�'!<<�����܈��U{�m%����֒�� d8�_����|(��3�6E��[�Z;�3�Ǡ��!�>g8�{�nPc�!��N�A�((E)�f��j�sGw��!T�<<H�Kkĉ^uB��7�-u� ��Kg}QvE��f���X|�s�(�-<���_ο�w��";(�Γ:���҂���M��e~�/�
��{������J�Q���:g�l�5h-P��xi輦~��F��f���,��#^����rYZ^��يF�<nP�+;N�E�\��"���@��A��=UÀ�[e��F�z�3�B�mB 4�`@�g�A�N|C�*���ĩ8��,-s��-�K��{��b���rnD4%�4��@0��|�^��ږ(��
-nY�,�3q��XZ�H��e~ځ��f!W�g-#�>
�p=5�{E���-�ӎ�e�Ұ��~��g\O��'9� �����_-|/t�F���[8�p�p��,������O�$�U�����ވ��0x8�F�t���ކ��^gY���kv��/�!��B�����Ӗ�v�[H��Ar�vnD�h�!E���E�#B�=K+E��y����zrT����<�^g�ۜ��M� �G�F#���FYێ����Hb!}Ή]ڡ��tfs�3��K����D�Q��J�ڐ��(,�@JG_9�r��"r6j������@�1�"� ����#ކA�)�PGצٲ�e$���XQ��+��b�E��r[�sO��9��>�=�yϹ�f�n��R���:f���g�A8�3����Ƨw���s#$3B�N�_���Ƭҹ+�O�W���@<��� �2�* &�u���UR�w˅��Ư��B��)"�I?%��g��{͊��y�sʂy�CB׬�OȲv�ID��c�aD�����R�O\Ԥb���W�6�����S�^���g�z�=���E�B�7�j���a^�R���0p���M�WlQV��*�K�?o�>��{��^�g�
Y�Z?����9g��Ա ����-ɏLH1��A�WZ]n�M�8�=�]��0h��Xh\��
��3|D@n�o���u)�jd�i�������R�O�!��t����Ъc!j���'�-�x�ʜ?z�ڏ�46;��|<�������p��;tE��p���t���f�_����nu̖���+��u�ަ�cs����z���9���T�0�V����<g;b��V[Ƹ|Y��6�a��QY�$��x Qev-m4�h�,�@�q����S7!5��g-�7�h���̸���dÌ�cxo���`��|�]K�R����º��g�
l��3<�+�Sf2+bhU�Q�4�zݤ��+�_��u��Z���R�a\1H�����"RC��~	�R����ٰ\������^O�&$+n� �Ld�b\�,\ i��)5�J_����ŤtJM����f����P�{�\o�R2t#�e��ܪӆ��\y�a��];9��g�PK   `��X�Y`�1u � /   images/d9bcf815-618f-4ab0-b416-9f611d86ef67.png�i8�o�7�$ɖ�$T�ʞ�[�R��,ٗ�lc�Zʖ6�	!;�ױ�,Cv3։�0��`0�巙��x^<o���⾎�a溮�<����9�y�HK������+�RP�VQP�=u��/��;����)��;�4�N�r��;W��߱������*Fz [���3
0,����������.	'w����廏���Ɵ��?9=9�Z�dl�l��ăR�-��c�/-k/�3x�Vt�k�4K
�1�V����JE3cx��\��E�݉�	5�����*,�Ђ]c;N'�Ȟ3�=IZHͽ���	U�qW��&��{Fܸ`��9s�'��%��s��J:+S�����*�&�5��^�0��������UR^���S�a��-��8��"�������ˍ��D:g��m�>@&�fJ`{�S��3��p�G,K�J.�����_p�0^�VmMQ�	Su�5���@y����?t���%���Y{^>5��z��~�ʕ8�Z��G7��fL���w&
��#Ks�R`��NLF^��n\~�z��D����S��w�66�-V�}��.+-�ۡO=S����	���u��|}O�Wڽ����QE&����Y��'\mJ/z`NSG�Y~`hK��Dn�V����m���4�[L*U�@>��à=hÃ��QJ�:vt���Gu�ƦP��X!��^��?�/?���S��D�S�y�:����}�jӨ���(=��z�n���kEb��[�������+�c�ς�5�#�-�F���6"\��~���/�䕸�����A��tM�?h��㗙��1�Y�h�;�B+Ч����G�����sycė��?|Q�c �0�n���è����q{5A�dk�s	�d�6k���Jd��f}`��9�;~�U��o��.pʊ��Mf�b*�Vm��^��{}��o�X[�[a�4#�BVMn�N��j�����t����:5��Enզ��ۮ�v�|�x,�&�Nٴ�����\s�)�<���"e�_%m�'�_�sń�[�\��B�7>�5�iP]����[�n4�X�4����_�|t3|�ӌ���]��70<�����`P;z��� ��h���� ����W.+�#C��������-b�:����.�=����]���[ ���]��#�7�����"�-��;)3�$�"W�������������ݩ�A1׀���fϱ��`�������ݶ�����uA�t���(lvޕ�?}�X}\熧J� K��5�ͅ���ȅ1e��Ȏ�>f׹�X)�����ɯ�>�7������鬛�֟���(c�FՂ��7������j��y��FD�br�fk�֚���d�M�9#9l/�nޮ�w�R)��Ctׯ0�:�L�dÓ�ݒ4v~ɂCތRG�Se�t֭:>W�u���-����՞d�v=�����ˇ�i}t{�J�8a���"����M)?kC98!M�͞��Hr{|sPG�q��[|7R��>R5�n$_%��6j�d���lGh;�@�5�em�ܞF?<Z'0������ڙ,���Ai>����yk�	jD_ƨ}���)S�ڮ�'��n��)	�7?t�~)k�m�X?uQ6�%>�׊��&�a��7���
G
��X�]v���iHmzJ�æ�ΘJԽ(w�\�j"�!���w�L֮���J�F[��JdA.�P}�.YZ�#����!��f�bf5�&���8��/	�3�|'3���5�.Li.%�c��4�%)�MB�-7�]o�L�,$�����U�n[���\�_')A�Y�u��E,'Ayq��@����ieH3�,�]J���֥<�d�`�ۓ(�l�<����ڏXo�aCkBZGƠ����}���w%q����Wfj�<$��q0*l����>��)P?KL�P��l��D��dh����;��.����x��є����B��<�hU;b:�;�Hl�����{��r���o4��+�M!nߞ=_p��h������/߉N�ňe�Y{�y,^$KҳCfl�p��7��Y\��>��^WC��O�2F<q3��;�8k|���TT�8��[9�>�oǮ���1u ���U��P��I�8Q2��z�V�G�s��\v=ܯ�lZ��u���aJ7N��<�'sUaܪ��3=ܯM��d0߀�1��0���E����a���:ı<��&P�?�C�Y�kL�ߧ}ث����
��"d0gVE����$ ���e��JK0pAl�aT���)�0��'�w�ssR^�ڦ�R�[x�P?�g���4{{Z��Ը]�҃���Ny�7����� �>��1�v���ޒ�Ĳ}YQW���=�V��I��|;_|� �o(u�$u�!�7ӃH�쮄M~P8D�P���f9�0�zp�^@�meE��V�/�Y]C����7�Օ�v�@Q7H��_y�BI���
r7�z�'#�lyca�S�JO���a���:7��Z/�&
3��Ż_&��~`ۗ���'qH�z1熹��������������ш�ܦ�̞x6�( �F+`���~n�Ѐ&:5�����~��������?���d��8�'�#67�)�wՀ�ٙ(���,*&��fr����ï�B�K+�����O�{B,R+G%��	�ݒ+u;̱����]y��5��e<�^���Z����.j�	��&ߩgו4Q����ky4���|9��_���렉���DB�~�j Qѷ�%YT/8Q�57��w������S#n#n��x�O`K����d��`���(	����|��;��n��A7�"Y(��'"M3�]o�G"���剢��z�y� Q�}n&AB�R1Q�,�XC�����kz�=A��B'��r��n�t<؞/5�C��ỊWfv�!{��E����[#��0j5��6f����
�1
��x�l��P������MT��i��_~4��������\EE�ʐ.?fZ�g��}��d���2M�J���픷*͉�>{q�	v&N�V�|�=�? 	1��R`h�ح-I@9�Oa��^?��/��0K��<(^0�{޸B����@�d�$�Ô�V�U�۸
د��E���Xd���w�"2�`k�vq8�㩚e_K��A*��/��Ar�^.U��T��V�g&�{�7����#5���7�I��'�u=��GU�׎'a4��fVy�hǐbv�l�� �:1	3�}�j�x-u�&���#�Jw� 8W�S�#&��>��2��.c;5�/~��Cv��������+�?���(�\b����Ts�_�,��f���� ��bO�DK^E����Jk�oq`�7ト����N���2���k`�$����iO�2��YC��26�\( �����{�}���I=;�������6#��W�7H���]���E`l��sĎ]*5��J�u� ����Sԅ۸F�S���пG�K�t�m1���L	��u9�� ���}�̯GI�]�(�jS�Eh��F��n	$$�ѫ6t�Z������v���?k�3�q�)}�?3��M��_\�
�p�``�>� ��k��<��c�7�&3�ր�r�R���rby�^c}e7-),��N�=�jA�-�����q}�|l;�厞{�Onї�� �	���|&_DF���K�4S Vݦ�LM�	���ӚYT�a��@o�ަT��d���T:�������uA~�ׅ�8P�L	���R�,��`a[�ǅI̱�X7�=<z>UP���h�.6��`�q%H���?5�}��by��,����q(�P\�_O6�\|����e-��L�(_`�AG	 �~�!3�FBNmӾ}�mV@(NQ���"��`OZ)	^�D6�?6 �Ca�˖G��$#��
�	cG���!*
vhԱ��gS
f����ܝ�d	Q�3Қ $q^�׎���T�N1�; ����Od��`�ٯR7��=/��B ��ǐ���Z�l9~��:�?���!~RG�)���vЇ=Zb�� ��X�����li�@3����
E�Ʊ%̇U���QWxS��"�Jj2%#�8�{Q�w2h��vG 3�'�1�E�jF�LF��VL�H�hEj,eʭ?J8]3�Re� 4����s�?u���w���ѡ�H�Y��Gd
���� Ay����ڸ��������u�<��2JH�|x�u)1CB,(; ���J%��o_�.6�åC�y��Ņ��
�鯴�a�7� "��0@�� Y/&g#q��S\L��UX��pP�9�ѫU!��7Ӎ@~/�Hg���ux���j���N�2�\�4��բQ#k@��`�����y�a��p��:�"Ã�Jg|@^	?��������#�gs��$�#,�v!=N�j8�I�������_�}��w1���=������е{:��9`y9>�,�^-U!̹ �G�(�$�8�l?_������Αqʰ�q��ݶ@�ˑ�_[�L�����sB*n�����F{4猸o����B���G,Uw���ŘU=W�%o�x�7�n��s%=�׉�#V���8�\bV�}��6ׇ����XMV1@�9Xau	��-79�՗FI���m �hߎk�n��þh�o���-8�z���;�w�㱔��p>󃎯���vW�%f~��?�	�ƺ��H���)�-��o^��vDk�0T�S�M��}���y>��eT�R�jH`�|��+���K{ќUj��0y ]$D�8v��j4���n}�$��^W#"}�Q����S�$��6nw ���Wu���V���6���m2k[�>�m���+:��JM��l�����S�@��bH"[P	��M��J��rD���x4l4I��M�\3��k��\6��,~�q��x�G����V<)�~�c�[7�p�;_f	dkY�jjD�Ǿ��Tr��Ԇ�h�Cdk�����P��y��7o�橎\R�2��%&�]�r�Р�\%����9PW���T7��F���2γ��Q�9S�Lɀ����0�!��̓������^�e�r���P����:�� v��׃�)�۳H7/��zޜ�V=��&!�r���ɳR��yO����VzdA>G�$�ߠo[!�$�$��;c��7�-k�����,	1;6��V~��_H��Z4w6u@�}ni�o�'�@�vQ/G/�`M<WT۵Z[��M��d
r���z�5���sN2?k���R0�����x3�0F)��2���i���l��g���햓(�ɍ�L���կ}+3��[���H�Vf� A�%Bvg�o��P٣@-k#��o�T�Z�;�@�N�h����b�ќ��+z�N-&K��&�3RJж�����+Pu����-�������k#�EYdr���LR_��Q�>#����Qk{vOG�}�1p�t}�G:���DC�;�����aZ���'y?�P���!p�I�I5oP=�?��T����gf�N&����s��� ��%Ę,��0%�U����=��QБ����&2K/8r(�X���:m���^�i�AK�Ҟے�VD��Y�<ih��L����-����^�4�î�X&��z���`b�I�a���7�@u1YR_���Y����a`��*� D~1�S7)!�U��dsa�ƿ��z����7hR���ҐA���	���kK���ai/_��e9�x�Z��@.!���.�@ϯ���b�Ҡō����6Pv�p2���������vB��i�����HI�T��U��I��'s��/�rgj�|�3�s���e���`�ܑ�p�"��o]�zU�T$���7�J�h�V9�&5:��|�iʐE�pGpL2�5�!ʱQ�rpL��zf�Z�N_4��T��&Q��Ɏ	CX$��fT���%<\��Hno��:���@h�=JJ�D���.`]�W�]џ`�S�HDJ���è��:g��p�Sw!�b�Ib�H��
B�H�tx�.z-�6�CmM����>Z���}��Z�d8� w�Dŕ4<q�~8��^��|��w�ގ(!|��oi�����h��O ����ȿ�E�)0sO��U+!���`�Ы�#�z��^PWWg���n���RƴvRs�������S��>�z��`,�M��d�]#�C�5[����F�5VOX�J~=���t�t0X��h�/c <yVұ�率S�z5D���y��<<���Rt��3-~:��/����{�w��z��FAd�5��E�����^g��IJ�H�-��ۮRddJx,-_Ơ=�Y�p:w�M6���r��Xl,q��,�wѣz��.�4~#�	3\�E���^*�#;O�ST(�PC�r�F��T M�� �l�di�=S�á����y�e�X������%$�������{F=��(">[�q������+�			�uaM�:�7s����$;�a�����Q3�N���?��#������
�ǿ��e���i��_	���wx�J���3��ƿĭ��o�ꑊNWLc[��d۷��w/��[�A!];� v��}Iz�Cnw������w���=´d�Rr-`ӆ$*Q8�*�/�C�u��۶O��˰p3b�&!ƣ��}8:�L�I>�;!���C{]!���~[bPN��_%֔�_
�W�<[��$-j��.��4_����;I⟄�$��b���3@��Yt?�>c�2{�;��4��T(�_�4
�{(���#VEWi
���8������l�/d%T���Բd�տX�*�ǩ�/�wMt�\�$
j��s�v>�'
���9:'.}�9{�7z�NP����P���!�%�?Nl����4�V�G��_����k|KѤ��H"�p�[T/�F��&	<�8V���;J��uu�==@q|&IC�ֳ���������裸���P��?��?b��,���=[u�[�$ӿIX�ʳ�%�7%p�84rZ�cyi���g����̦��~���d�Mx��%���(8�����BJ`���� �Gw��ɨ] ��֜�!q�Rq�#Gl�%Fn�D��Ld�l��J������I���57rVY�t�t��AM�Jѓ*e�����:'ٮK��|c���Eຟ�6f��[T�LIم>���{Ù��ʑf{��L��٣�n���4�*������h�1&W[kg�j0���Ay�lz�EAU��WjްAM�#�=��<Z�j�]��Zs������_m��'�W�?_йa�g^��!�dj�S�g5��v��V��2�[����L(�j�8'*�ش
�	l3�	��ڕ�녵Q�I���g���!�S�Q���h�k'e_/�j����^s=�X��"og	��"L@V.�	]l��bU>�K����c�5?Q�X�e���9h��rt��8]��u?JW�]�9�����zE�e�_pή0*�nQZ�q5�^��&�����T@�eo�7�a*&��)�.�v�\���A7��[�FZἌ�����B�r�D]Z�Z���V���~8s_��6���7Q��	�\?C�s�'E�n�M~�1B��ؒ�_�V��2��E�~Q�?%ǅ������#Mڌ�Ka���0<!��/<GH���;Ұ�P��y鄤ǭ ��{������D�~U#�U����N��}�hAQ�6*
ݞ�
d��� |4��G#��n��hY3U{Y�B͐XG8�
g#�����l j�����#X�P�G*�H�V��eu����A��vO��0,%~\����r�L�������{1WU5�߱�M�,���N^�C-�:k�qmο���aJQ����r�
uo��q*�B�9���p�ψ����E�O	���A���4o���TW4��8Z`=�)Yv��An��J��á�漣mE�d7@n��s�/���u"�}�5G&�Z�,[�����/��Qv�y3vx�s�Kxm����1����ߣ�G=�������HM�D~K�1_�
�ҎxU&u?J2F3䩝B�>apw�u�E^nbV3?����l\�A�O����M�����d�~Mq�R=J�CZȑ��<�䍭�Ŏ���A�a.W��)�4����I�3�PS�4O�~��o��W�>�y��z�z0�OP�F'R?��h�>�:��j��I�|{���ds��JB�
�RX��}�Qڑ�|������a,�3��m��+�w����������"#,d�/&�����=�3���u��/LZ>D�1
L:4g��d]��hBx��m��h����nyjb�l_<+J8�o?2�F�h�����!qZ��08��v� ����q��/�������o;�55�}$i����^Z�b�ъ���[�Æݮ5����/N���)%s���N@��|˄L��:Iƪ�M'��
W�Ogv#���)�3zBw��@7���οpm����w�N�z5�Rچ����G��VT���:0���*�2�����c��/�8�::�4��e*���v��ێFÈ��2�[l�~Q���1�E:���ԌS���Y� Kg7>oܭ�g�q>�3rۖ�40��Ƌ�h�W]�1�{��j\4!�͸��~�H}�3�$���"�լ��W �A�\|�Y�<ٮ��� ��bÿ+���\ܐ���7Ӡ�X޸~+��`9d�-���w^T�y�cA¬��m�w��ܜ���_�cż��aT�/��$�"mB�j�=�	m9�یC�	��c(QC�5;�z�3H���A������y���[� B��SY�"#��c��)�Н&��ٷ�v	��j0���2�<l���ug�=AuMt�)f��{ϙ��^W���3��p{�r��ɸ_��7G���%���ϏiKtV�d9�
S���vy���]���D4*2N��JI&��[���?5c�����B�j�U�� ��넜E�O��B��r���^网И{MM�xS��u�'v�+$eΪZ��(R�v�z.!���<`����t|�W��Q�*��K�q����_�q3��<�V":6�2zuۧ����^�u���*��z���uJU<��'�v'��;~��
��������
�ͪ��Q#�2�#{�cJ��L�^�����"�����u^�����$���K�a1���iY�Sn�IR�[�������\Nw�l����S�p(��9r)t��j
�:p��o<�7GdS���l]���ud�S��G�c� ����ƃ�%b�Qp���?΂2ow'��p8���)y��� ��� ��s,-ȇ��l�@��[EvYΡ����[j�*{�␢~��t�q���m��q�S�v��n�T�1��׮o�" 5�Ef2Տ� �|�z�GF�q��e˻_�d^D�xPƮp�4e1�y	�W!1���o�g�v�ض�)>����r���{��x�.@��g�=+Q�8S�@��H��֕m_�߬U�I��|��*�G)����Vg��͏�R{w��]��q|ٍr��M���	K<�W�~B�	����p���Pq𰁊�ʫ���7�&��_�dZh���	^�)�T��o����1�S��-�N���Lo���4��ZZ?��}�C.Q������Ml�;F �lT�Q.��{�e�L6G��4P뢍{��'��rVk�~�g�u7F�7y�e���9��JZ�R;Lz9�1��wOe>6ջ�?�V5#ZM��w�jAG�����\K�@�����"�n�*���������'�t�o)�8y;(�??�Fm$�u������^�r�s#��U���ә�U������)e��Sg)��N�9z���A����]���S�]S�ِ�Kx���.3$9�`q0���5=�Ҵ܈^��ے�ǟFm�X�Y���8%����#m"�?p�b(��)�<��/��ɖ�FD���3�}��|X*N�%�Ѻ +��hQ���b��h�����!�Q���h���j*�N�,����%�+��{:O�)���4�T�"����FύSQ^,�-��S�mŅ�E�4N��&q,k}.�`F[�)����,���DnS�gE��U��t�a����)�g0\A2EC2:�0�Ы���9�{c�$�7pV�W�yZ��Y4[c�i	�}��YO�5��\��	���|�g]��[�ygy�I�aaH���2�З7Df������!L>w�W7ey�N�Y�u�k}s����5��׈������9S�K�����}GZ�i�T����Em�)�㳫���g�1��J�����3$�yTk����S�,d!4����2�J+�|��KW��6��V;��a ���P���&W�
���ǫf���#�!)M���0#' ���)��߆"���k �`�D ���`���mR�����	��������2c^����]�;��G���^���e�4(����C��m���XZHē�W�_|��;wQ�^�Ԁޘ��rԷF�3���[,��@�CBI�9��$���Z��Er�<��#�1a�ء�ຜ`#��xX#�e\a��˻�u��1�S`���3��b��C�/o�S�G�esY �&�$;դ��Q�{�;,��I������8Iėʋ`ռ��1���&+c"^��!}>F��N��=��X%hx���������!x�;?�[Yo���%.Z�휤�%���G�i�7�6�ؠk����rx��	��Sd�U�9=����RX-o#.��1hA��[�z���VS�(ٱG�aߪ"�~�p�*�U�����8y�9�
}P�҇6ұM��"��x���3��u�g��#m���Þ��
�d�a��6��g�\����f�{��*R�I���nl7�b}=*���c];`o�W��GF�Bc�toZa�PEeiڅ=�S�$Զ$C|e,^	��M-�iɃ��M<�V������Q�W�b���;Uz�e�Ӱ|�r���������t�*��r���5���&�{g��r����m3��Y� ����	v		�(�i�c�k�m�����e�T�$C��KQ�l>�.�l�Z v�M肇����eV(`�M������/��!�2ϔ�9b>2��T�n;�^Ξ�����X���z�c�6w:�ADH�<闟{�qI��A� *�Л���6U
?��M�L�) pʾ$�>�D��I!�1�_�ޖ�-�h�3�v��s��^�qǣ��M��G����,�X��$nW`��9Im�(�R�~���L���q�j�����m���=ыݥ�蠻���l���̛7V(�7��NB��Ch��s�3�= ��M� ��ۈqO�Fp�$,p}��ru�8��4K,S�q�:ka�	N�o��)��w��W�k���'c)�>��i�!ۭ�V=����<��f�}<f1�4���,����� ��sR��j�3[�<��`Eϊh�����XZd�!��Y%8o�z*�C�Cn� B,�G���cF��`N �6���l6����9dɊ��������� 1�ŀ
�EOZ0@L�B#�=@@��t���5 �P�pƯ|�N!ʲ��y,�OӠU���,�rK�R�E�25˯��Zze�HU4<jܭE�=��gX'�0.$����ܤ>�;{+X�ޝK��!M���T�LV]����B�����xȜX�a՛4w~e������&���m���ԋ���+���e5T��&�o<z�^����iG�^�H����<�U�Q���p���p"��cv��v/��YV�[�B *^-�tW]�Uy��5�vR�Y�H�V�@B�5��%�zN��Wt3`���RD�5��HD����.���[ ��M�l�#�n/���"H4)ؾ&��gC�M��6�k:L�M� _YU�4������l��Q������vے��\�������ӎw��A��+���n0Yq*���Is�l�&j*����w��$��O�:�6����ɪ˽"z7o�U�4�aO�?��>{S����r�#%�[Eme���%.C,��`2�G=�W��D����(I�([�Z`L��2g�@d�|��v5��ث{�2=C,ף�ԆGW�Foz�s 9M��HsT����Ve��`�i7�D�#6}�~��~vRy|"��5 ꠦZ�K{��3Bt�%L��3�5n&����"��?۩��1↋s������Iޏ.W�X�< {3d�#�ﳠZ�k2��AF��Tmp��6)hqa�v�vT��X��abi:���ߣrn����R�@б�^G���tV��a��Y)m�:����H��Io;X��:�x���q��N��8�P�p6}��w�+i�O޺[^�ѓ��>�.�~��j�rNt�t2�L�����ߥ�z���n��c��H(�(�W=DrhUiR
}V���ػ�?4�sr��͗�,D|4���3�Z��Զz��z����M�2uӲL%{Yd�:���k�,V�86T�����=cצ�X�/M��+������!5�XW�s yIt�w5f����ޤ#�f��m�B?��d[�������~ztm��Hj!��)���`]e׎�����]�6s;��[o=�+�ACM5�[��+R{�P�d.UL�3}-�V� �+���5%�� c���̆Ӗ��[ �!n�7J$&35�������L�ޏ��	hҊ����<
\壢f����q��'�NJ�#��e�Nk��!n�O��.#:��-��~�iO�0�j>rw�
�M.�.#v��l�����¢��h�85���%�!bR�{|3���ڡ;i�I_�UGO�C���� ����-�j�a"�G�Ku#P?c*����P�G���5�~���1~*���uP���q�x�P�2��N���{��-��\uq��#�헱�~sQp��<��* � f+���#�\��Pi���-pX}������=c;	!E���-��ћ,�C�#��#n�gD��S��c�Y��ԯ��V}���GH}����p�����>�?�t��ҦgY����U�H]�ˆ[~V�B�_c�t�ռ��K��if�N+;l�e�����齢�����AH�$!B�gȭ&v֣�K��#wkX;I���H�]����<4��[8�>݃{�P����v��+�as�g/2��O0����y��&��m+6��f�y���Ue������iy?��MX��RN�\#k%^dۡc���ٚ���{�u��t��:�b4^��
�/m?��S"�E�RQ�%��"{NH,�f����~�u������s�������&����j$�)]�D��(��W��6 A��%�%*!'h�0m��GWI��i:g;��ݐ�Ac�"��2����J:�u"�"����-���4�/����Ռ� ��x5s�D�{��N�E'��6�O������k~��F��k4�0mYXZ�A�N�5u�v��-+/@�I�8f��4�j9�[d�^׳Q��.�G�,y��8
;2����#���C���C`��<�h�\���q2��G�o��aZ���״��,�1����-�V8�&�W�\}����*f� �qDL��8�{ԛ&�<> ��0�#��%F�d� u/��AN�7R�WA	=��svħ���O'c��[����cX(�{�gh:Ԝ~�ǹ�0=�z��?�ּ��pF�bM��*�_�Y*����t-�0�(J�G�4���(c�QI��G1\�\����}q1���#t��X�σ�N�;`_��9)�ꓰcOla q��D<����L�(��$��.�Sb�����4 )�����i>�k?JV7�\�|�&�+�0��/�F�k�}~ͤ���F����H�Dg�m�"�����
�a=��K�����S���v��������5d[ڕ��Uiϭ1nT^NV)�t�c=��K� VXm��=���cȂ����e��x������hE[�q��9�t�5Σz������Z�ߒ?�rp0���������QΆi�,8(�2�9�\R�_�*,�x�i(ԝm٭��On�eo��j\�S�u�)����󺌾��k��s�h�~MZ���4��C�;s��N�Gԯ�ҏD��T�$ܻPƛ.��8��4i��I����o��nq�l2QG��F+�b�u��O��-1��6u��Ptv+l8��P�Hs��}�J���H��)�BφԳf؄n�L'�����ޫRp�V�].�Z���4��G��Dߏ����hs�=�ͽ$�%�-.0�������{�1k�S]����#s*1��֘��GBG)�,���_���9�0��ʠv�q/7g�[��,�@e~)�𙓾zT�f$�\�V�ǌI�-�k�E	�X��X��� �iC���c�lSB[���)E|<~��"�B��@)@k[8��p��KO�I���cƗ�J���m�~O�tq��W`�ײ��2/Z�؄��^!��.<�dm�1��\�Q�G���Lok98���M* +k�E�� Z�[
��dԴ;���;*�H�T.aʲ�4�::԰(Y+c��8���$	U{�U�����FH�4��gjTֹ��>���M��y+�U�֋;�e^�����y�Eq�$�sfrv���������A�6=CL6�;�+�y/Y|$�Cok�t"\i-�1>o.?=�`>G�G�)�q�-��z�sC�m߇��~�;�G �c4EP\�un�薧L��$��*C�3x��K�c�K�CP�߳�^�'۪��[��Z���|��k����N�E����XPHSmڨY�A��s�&j����~睉]�*���Bf[�e��w�nG�[��i��5Y�K��p�r�}��'�H�P������G���O��qx>=	?m�eX��z���a����57�`�=��7�R�	�q'̟����49�*Q8�q�Jw���&~�4y�(3S�C��+z #�e9NО^jQ;:L��	7T�m��̡i����D>J�d��L�o�ߩ������`ϕg�Y5a�6z�G��DWۧr�	z�:�R�-G5��E/!���ٞ-Ê��l'�m+��,��Z����L�T&�c6��[r��K��C����c0����6�Ǻ�.���.p�f�p^>^�X'a���L �L�5~m�ԋ�V@6�O6�xwZ�e؎�͇����>?�>��*�@���*H��0l��-�B�B"�o�7����cA���jk����/��v��7��*���w,�l�A�Pa�A�ϓ�!���I�� �������%j�{����j��`xLsj7��d�gA��|�t�\,��t�}��N'�[AhH�X�N� �X�6Sx��)��О���^�6�š�H��œQ�`�%i�"l^]A���������wj�l~ւ|�����I����ߊ^[{��I��l%j�b�W��K��7��!���!��d"�?� �?����o?�L��&��:wZŗ��{v�s\̨�N&q�@;�t��M"�ӵj���_���|G`d^jWVq voT������<���.��p������;SdԱ�T�^�Q�h�*x*Y^� �͉�5�b���	��������%fs#��l(SO=�3=�D}ϗ�n�o�����qc�g2��e�M�.�[~�
�_���RV��~�ih�2b�����m?��>��}4	�~��w�D��Tz<�H�uP�O��� 
��8T��k�pix&}���J�rK%�>F{~��H�_C��X}��-S���W(�x��Ąn��W:Q﫾�+M�����`OU���k+�rߞR����^�2"y�,����j��G:Ѓ6^���.u���r���x�ڢ,
�����2gw%֡���I�`!��RX����l�y���9-��̎��-�8
4[�K��	E��n�a�U�+O$=�Ͻ!K�'JS�]����<�b�A�nq��ې�C-��d���ġ'c�/5���ŏ��#Ó���S����m<�m�B	�FT`��۞:�"`W��$���߁zS�W=�f��F%̲�;����6|.�砛��.�]%
I�l� 5��d,�}pK4}٩�]�3��s*m"��ؠ���ۈ6��	d�������_Go��˜=y۵!�Nue\�*�!�2_#i���S���W����1F  ɣ#�ج��e���� !���G��� ��Z6Ѯ�>���*�<�r�' ~K*҉Aq�i]�X<��>*uO�
������ӏ�׵޷p'2�d�`\ev�d����l�nk*��2���0�$��M~1��1�U��?D�ΛZ�zKa��)9�\�R��>�6J:J�Q}ݻ�{W�ߟ}��E�D�9���2���v��d���FAU�U����b�j��ڸx�|d����Qq��.�%�*�N	{�Bl$p�\ש:�v'-i��U�y9�B���"�:>8}jp�����< i�#O�Z�5��u�5��STsBOk�/ii�V��~(��*�.~
���ڵ���'�E��K�f� ����Լ��A�(�X�L2��UE�"�<bam�Zv܋ӳ(�'j���M~ԕ�7K�a���`����cOa���W�rs-�-h��L���rAo9��*��i/��m��������Ο��*�`4��B�9!C�PH�%�7���_pY��/x�$�J��\ot~���_�2�ypR�UL�شnޛ7өV�a��<�ٰƎ�w[gec� �Y-����N�t��M���[�/m-f)EmN^��J���~��"ǁD���qi�ril��$yZ�9�~�؝,�/?X�U��♳6SI����;и�����G9�|/���w�DA�)Აj�F��K�K���u(��蓠S����������rY,nv�����ΐ{
�R������3da�Ud�$$�ҝ�r�ժn`K��bc�mv*���ߊ�Ka�eiS���N���k�17��
�W�R��s3�؟N)͏���/���|��Y�p�2[L��lJ]�i�e�p��R=���B�s��^B_i�٤��N������{���'2�m�|̔}n���TK��|��!�^]Y�#� 92�wS��Mfm�=b�o��沸0�M� ���l{���͜$c�茁h\�)���d��f+�ـ�W���'9�R��R�2�0�m�o�=u�H� `I��E��R�v �c�bn��L�l�W{���(Ȁ���~�)��9J+a���@p���R��y��O'����	c:�~��Ol�a)5="䍿h�W�����l���غ갨��� ��J�tw���
H))-�]K.-!",�)��ݱ��tw�K/��<��������3sf�=3��s��D!�m���O�ZW7���E�*�}�;m�т4������.�,�S�F�m/[�P��YmM��\j��yxrZ����5�m4��7E~Z��v�-�92���}uO�k~�)B�O}%�^���^��{��!x�9189��Z$��Z"�{��R��<D�^X�]%@.�=4�Z;��,Q�Z�D�'�ĕ����Dx
�D���p�ʹ�q;��'�a�1ۍ�ӕ�'�[��y�bY��*H��%<	�Z.=��$ΐ/{�ɯ��ܘ���𑆫wC�DO�$�弣o���FK`ȴ=3{�G��킽�^՗�^:������ݙ;T�6��mϷ�tR�E4�/�^;�=�:,^7w��O_�W�5;�����[��T,�T���HLT�Υ?��-~J6����[AL�r��:-�+�zN�
�%G�Y�f����� ?p��Xdc�P��~�a���\�-��ܓMT�M�o���G>6K������%`�;��{��;�P�U�������l�y6Nܜ-���W?E!Y�j�6t�M��ƍ�1��� *J��
^�c�*^���??���PV��,{y��7���;qu�(6�.�@Q9���g�<d�׻G&Z̋�1Fev7����y������b�9-c.��Xya�y;;����̯oiֶ���r<{H�{r�	�Nf�)j��\L�[ �L'�#ƌ�@��g_V� �r-fl-9/�LU��	b!�`qq�K�~��Jdk�h�V��~cc�e���Ԣ�k_!�����Łg���֧a$�l�[��۞�0b-�l���F�e�s����b��蕚�G�u��z~�Y&䵈6ŏ��eXb"�a�Z?��&�RS�.�̞��ü	'm����݅@p�l��V�ڒ����~��5�p8�y�O��)��o�4;P�N�r�%��=�:�Ĩ�Mk-����о&S��2�l���@RzX��Ր�J$����k���ރ��Y�}ө[0%��iO|z�;�N$��E3=&�U��4)ꭏ��&WWZW��n��[�����K�..�;9l���AΔ(�~o���E�_���QCTc�����`X^���z~i��
�(ew��p=��^ȶx<��C�^w���]���Z�5_���ߋ�]�ὒ�~�����ݸi���q���>����W��r|*�t��c�nލ�kQә�HilJv�e�6��`h`W��N8� �V8K������s�j`����@�����@�tK'�.J��Ծ'/(�\�<�w��iyb�#wrΝ���ij��WV{3���)]7~�Mo�:�N�M"_�@��݀ы��۫�d���i6��Tf�Ļ�P�m�&��mE�ĭV���8�i����H11��$����ҋA�Z����gv��g���W�ơ�({��G����ͧt��(�Z���X��X��#5n/GK�����%��غ���掮�CG�[X=(��?[�KNW'E����x��y���.���Ɠ�,t�z~�\�8�+&ى������g��pG^��7&7����J�q���oO�zؠ�]_�V�c��B�$��0n�ٸ9&\y��>����<�4P��؛{�^ �z[��pa��xYz������V00O����/Hd��@t�n)���@A�:}�k�2uq5{��?Ax{M��s�>����floB����^]W�nu]E��&���JS���`��M@b��5^�|�<���g�����2�`x�bS��X8�3��B �3�q���F�U/+�D���.E�9ԍg(��q��
�8�6g���`H���V{]�9�p�j��� ��*P6�:=>2�५)j��4�̓�Y>�7�H��4$p��e���������e]܅M��M�@�T��˦��ů��E�<Ay.�	����W�+K�}�d�<Uz���K�G��n�T�BS:�V�z��fH�n��#��ܐ����=*4����[_{v|}�u���kQ��h{߽�F֥��Y�:ps|Q�^����LP�_Z�6���O�D`�{��Ⱥ����Vh����l�D����J�.<rW�g��ڇ��\#��Yw�b�A�����Z��1Z�l�g��S*��YBkj�wI�|����T���jٶ���^��͜ΰ�u��ċEG�#��$-9��ܫ�����.����o�`}I�[�ZoA��ו���T�x�s=���S������96�D������/%�����6~�6f�خ�_̻*AZ�V)��J�zy3p��%gYX^��mf�����O4,�}3�i�!�yq� �ڍ�P½uN��0,0���"٧�{`��AR]�Y�]�O���
O\�H�y��A�����Bh
���8Y�^����`��S����B�׾��`̀J�D�M��#Ђ<F��ނy^����s����.Qffo�ԍg
���\ΐ�R�������P�)���D���)X;6g��k<��� ��d���eer/o�7ٕ��t�������%�d�Igy��������i�(+�XLκ��1����ucq�2;�xC�Ş천��8q������/�+�?�u��uYvv��λu�OO5�n,�컻0�s����ܔD�^� �"�.Y��I�bt�E�����/Pw�ش�`�;UHD���݄j�� ����t�S�v���-}_v�ؚ9Pt�S��f���e_T=��&�2��I��4wUD�0/�E�j�\�z�0�ۛC���|â��_}�q��ƛ���b����Ƨ�=���F��5�=8���<M�����j����y�	M��Pu�������0��:��D׭)���-#xBA�/���Y�#����\�1�I�A����q�������c*!r9ֈ�-���t+ʍ83�m�̈́�:AJ_r�M���k��oOҔ�'��L��V3Wה=}1zs�A�V/%NzCm��gka���<��A�w� ��ᴹXН����aS���x�������ݶ��YuZl�V`3����=#*|d���p��_N^!~j�{��Ԕ{��|ih�K��c*Z<\�q����-N���Z���@�p���(�xiq���o�@T	`�%��x$*�|�B��J��v�":l':B��U+X~�(���:'����͕���>�,�^����X�MK��`�'{�X��(0\��s��v8�ڒ�8�}h��昼8˱[Y�}lP�=��	$bz
5Y�N8S�6�d��k�_����f��j�s>��U�p���ɰ>Z���E�o��ދ��d}[�-�[�Ѽ���@�'����9v���/�@ݏ^x��A`xj-� U��[��h�*P��^�� �aBV�-P�Խh�֠��Jrz�	U~CU���섁��G�	ۅ ��=0is�_�[22�E��'�}�@�µn�lh�X��Ȳ�*���[h	��Юx~���&�o�$U�;�}�WN���L���{X���E��C{0���،1m
z���d$�%��=�U�%f�E����#��j_�<���5r򥥔[7�K��IOe(QWU��%���?�nk��V�}��;$E���r|�?���~��r�|��z�e<��D��AIh�-CA��xp�*��"��NWC�u�7�*��<�	�v�8'��D��	�=i/��{L^gsS���.k�'[��L���x�&�ʉ��U�?��X����g��]�r\�tx����c6�xOuCp���@��3}m��m���� D�ۡܻ��P>���&�X��;̺�^���x�����ȇ9����S�$K�]ag����u�Ea���q"��JcD��#�/>���s���!���!�f�ê�K�\��9΀�ڄ~�vr�܌o�`���u�S�	r���_G��Ԟ�gN`#K{L�Z����^y��|}�I�j�}
81U��.�:[��%����2o�t2E_�r�?f��{ZN?�;�B��}A�޴����Y�?��e��/�i0S�'��݈��O9�ܵ��%4H���|������+���o'"J�6���L�����>�����gJ��r���	�	l�����P?�,��:q�>�ae�ϧ�b�Q�:0�5Ȯ{�p����|��DS��܃zFfXZ��D}��HQV��V"ӣ��7�̧���\L	��mkO�b%\�*|�T�cp`ꨄCd��额���YH��f�c]��'��iE�D@~�y:a�?�����滼�f[m���U9��'y��t�|Vl���G��a����O�?����F�|�>O���&�9��W
UV?+�l�_��:V7��^����hN��v��
��/CE�:8J��qUw���8o�~�z����"+1�w+��pKz���_���7FC��#�����	^N�ӐNN��B��!��j�|�V�o�?��GuNb�<eg�b�X��4D���A@@�C:��4b]ޫ췇2������헚��s�����TCm��Yr`|�B��؍��kT�I�@}2�=��o>�8�d���Ha�]� �;y����S�;�,t�� R����^��o<����g�G�Q�6��,>,��V�'4�y�B��h�M�r���
�C��Cx?&+u�A(le����^��FJ�viН]3���A�8�h�0�T=�p��X@���K0.@��H7_�*?��?����s�g�U�68i�����a.�y�� M9��L��@���F�&�!���~��[�b���/�O�HZ��>�po�s�a�1����w��=�B�'Ц֣���]��q�E��Qq��:�u'����/�C���6�������ޠ�/��YNn�xgǷ�!�j�	�ѳ
���/4R%�?�'��nn�JGg��<�h`+�Ɨ�߅���}�����KF�']qm�1-ܗ��7t>L!���.|p$g�����L�(�a�4�騥E������~z��$W_���w�nY�켹u�����Y<BR�����l��:���˥/�p=��F?�X�B���}�j�wJ5�w���f�:;�.�3��0O��,��	Z��]�ɠ���u�V%��_�s��X=�		�9 j �/��5*⹍lV�L���5�TX/���3B���l!x��t-.E~���ܒ�	4G�q�6��*@;
q�Z4M�?��jy��߉ rs�b|rD�]��`�guM�GUhX�C��Aa: ��1�_�J��k��W�J�8�k8&�'EQmۣ�	;����V�S�F���/�(�[2��o6��ԋx�2��C<��b������i��lÿ�>ӓ	t��D�7��^$$��^�m'�������g;8Ʉv!�Τ�b9�Q����V��γ���7��ez�$a�8ߗ�2��dj��w,Ӳ��l�]��Yu���c�*���'�Aٞ����ੌ�(���z'*@�N�hu��teZ�>k��hjɪE6��@�]��dĬ��������8��@-�U]��e�0��V�1ѧKo�)�Q=����d�,2���l2�@]���

�߯,�91�������2� 6�lg�:��gPږ��v���e�>_���m��o˭��0�G��N}�s�F����������a����W�LUq�~���4�������>Y���A�m�����ζ���Bw�;Ӯ�@��dm��������c�r�[�ӮIU�A#�=�*O7�cΣ�Ku���+���c�7�<�{�(M��.��7ݷ�_q�^��a}{�<ʓ�n�˰���i������K�*wD��Ϲ'�9�~�lLw��&z�Z�D]��o?F�)谄�"N�������G4_3�@P��>P-@6Rj]���S��EͲr��NK�2te�n oQ�\��%н��ʩiyPJ�����FSs���*�t�owI��&i2L@W�b�X����4��jz`�4���Xj��rҾ��r�hx�1A#򰼡<�.U%M-�O�L���6o����pѐ��M7���\�|�;
�n�C�^(S�RN��`�P��y��Ki��4j^f#A��_O�.;U, �͂��Z�p#<8:b|���
�Aw�ݸ)���G�QF�6��x������ #����P#��Ȓ��R���Z����r�Z�;�1�b
.�����_]�O���j'�JY�W6��|4���q1�ò�
��"ɡ�_|AXXw5U�9����{��)�-��(8�K��9(5�H�	f����d�-c0��\���R7��1��k��*�P��)^��󛾰Ǥ2͔,`_�C� T�f�^ x[m��k+��4��eΤ���Pͻ!��@/@-�]�9*�4C0z�us�A��>���h�40�=�g̴3��2hP���=-n����]J�C���2��͵�.�~��l+3X<����j�2Y������C_e*4K8�WGʹƤG��r_���+�$�	
+O;	��:k�we��	B=�{�(�^��`!ĩ6�D)��[�Hq��lx_�?��.���M�6�28>;�4Ң�ұ�5W�����?R�?��c����p�,�7��G�g������5����u:�z��b �T{%*f��X��9>�X!g�"�@E�B�K����Ҫq-F%���1�L^@<�lz>y>�s����xL��,)�Wڼ֧]�;+v���K�����U�CU��R+�����d<�x�H��w��w�����V��m��kmqS������=��x͂$ˋ7;�ʲ���i��K����:��G�]���T3�l�b�">,u��ǥ!fM��E��(X�itIq��. ��N���C��DΖ�z�X���U�*%��0�M��ۘV�|r�z��a{sԉ�\������n���b���C�����af��3�:�� �^��+2ĚO)""���7<�(���>�+%$%:;�[God�oS���ؗ�%�q��!�sԣ�U3V\��1���\�0��A���1V�4b�*���>O*��ׇcv��ZOE.���ɡ�\���K�mk0�q��s��l�M}��T�߈��Y_�+P����ͭ�+0�8|�CV	ׇ\7dԷW\,��C��^8�ɩ��I
��ݙ�c��\�1��9���)ݢ�*Vđȶ��0ry���w��jN?R>��#)D;��;sXP�I�̈́��?���V@���K�[L�b��Yj��@��:)ȿ
�K� �M�O���~[���榊��g���=a�;�.��wP���}/��@��9E��g]��A��S]?�͑�O_��Ƿ���u�̷~�1�y�h�b~���M}��<�5�$zə[ȯ1�k ���V��>l:�&�nS�8Z.?Zߠ��ku_t�i�L��ۓ�ڠ�ߧ?;y�L��5�`������s#8/�p>q8Tq�J�q_�k�;�>�^�A�{�{k+����Z4y���|�S>��pnLf��i�,�������1� �����o7��*�+yP��!���,K�M�v�4�N�sL���vo�5�و��Η���D���Z^�G�ܽ�:�j���ȱ��t!����~�(=!9;�ߧn3W�!^1+���L���6�0Bح�,������@f� `Ӕ���?1	��K+�!����WRݢE�m{�����^���o�cD3Dh�֎�Gz�����~����P�9�1�j�z:U&1[)h]=�b��H�������!��A�If��4��8E�1U��P���V�J'��?�f��+�%���~���<���fV��s�0�C]5��a��A@q����:O��~�*��H2�R��C�\f1T�>�x`H"�9�qQ7O�j�j��K���yz\l��f��B�����8���~v�TMmB��u����͔f��;�:��Y����N|>�)f�ZJ�_���vx���35;�*+p���'\W��j�����-ؖ�L��b�z���p�$��C|@)�+kq�
�L��Jη)�i���I1�o�E<����8�q����xڜfc#d�ߵ��#,�h��k��R#�L'7����<��7���$���c����FQ�����u�3X�@��ό���*u{%��a0?r����	K��
��b�w$w�X��x\���I�$�)����������Ι�3>��g!�2fs�������(��	Mg�;P�_@�V�ܯ�d�_d�L*��ڹ��|U�o���{��b�P����虹e�����q����~Ɩ�@#&��Ѣ�e���_�;��"��ݓeޡ��Y�x��r6@k��r+؃���ˆ�J!�
R�0��ϓ���oi���G8��7��	�N�7�1�0:�q����w�̉J���|m� @|�_,P�ϗ���B��������`����3m-�4j��j��R���ȓY>���c#F��ȴNYl�Q��$��WV)ǣ�Z�_�B{z�̭���'	��9�h&�4x���.����@��i.��B�3�(u�h6��Sʿ�������@qW,nBy��E�����; ��{����V����3[d/rЧtzc0�,%�k���e���:祾����I�#���P��zr'��3����rX!,�+e��hEw�д��������1�׃��z�K���U��Y@,b�Sr������u�YHA����Qc�dF?1�[������q��hJ�^B6�q�X'�屛��E�rm���{8E눯�����'$c�0A��h��y�7z���P*�k�'��!
���XW	<5j�!'t�t=�i�9�Kv�F%b~s��/|#ھ��a��߲�tU���j+jX*�df���?��)t���)� (�Ťdw�,.���Yz�w��?��_Gp��߯Ь�-�a8����%���X�Uǡ��lz'�3������f\U!V�7a��,qIհq)؜���\��1��r(|�4�x��o��p:������ٚ7�}��������{��x�+��QsD6�L�iZUk��FH+��QW�#��;AU����Æ��������)�`��  2��?.���X�+�����\%Y�@���$I���Z����-�,^Xt��e̿�tg �d�g��>7J�)���c�᎕;% �lA랝�j���n��d飷f��t�^h5�f�a&.�0W*��d�el'��Z�dW�-�靽h��Y!����j8J�Q����Lf�`u��jz�9���ͧ��lt�ɤ�@�ӥ��4��PS���2�oy���J�b�����]����V2~wۨ.�N��Tewh�+�2�d��W��5�q�7�Ȉ���]�K�,:��o��/�G�Rί����q�ϯ�=�z�U�2>�z��;�wo��1�(�`�{/�rG2�;WAcB�>�;W�Jq:cG�&W5X���$�?z�a����P��N�����ӫpC}��LG��*��q�M��7���Zī�>��J��<r��E�p^.������@<���-
�x�覈@+O���Y1�ٶ��9<t^P���k�`=���5G��ͣ=xծ���Y��Ge�!πd6#�7��V���X;�dCG�v��S�H�A�Q׵-h���S���B#�e�q\����WQ׳�^���w 4_Z����I����,�_�5륞�+|�b#��WC�$?ų���_�������L�<�PW{�;b����]������vA�Խ�/J4���K}�?�axdw�g,��y���:ٳY�ܑ	�/�����p���E�^y�D�p�S��ϲj��ߩʛ7E���[|QDwm��!�,?�b����?��'��g9>Hl�H&��~f{A+��΢xY=�&W��im)��'8��m��up�03�g��O	���"��_�`���S1r4����C*VR")#@��*T�?wJ�1;��g���7��A��ʏ.����L�E�C�f�F&����,\���j6��\W��
��h��#��Q�?1[�kF�Rt�%d�\�3��$�R����gt��F���=��O8K�aEE�5"g��ۦX�bh �5K�Y)���5��zx����9Z�0PG��$�ٽv2�>̾�J��ٱJط�N;X�2)���9t� �ϗ����_���8d5C^����(�K�%K�$�F��L�'ۍC+E��	����WA�Nu��5a � �֝�ϗ�o�I�2�(�*Ә� ;ag͐z*6'b�+��Gu[�x�;����BG�u��'\��F���6�dȼTG�����`���w�<��e��8���́|��{t��2:i3-'eI�a���c^G��͏!� k�*r�!B�Y
��P6r���I��H������a��Z[�X�"����JQ�shG��oQ{_�u�1̃\���&���;���8��@O8-��`���QJ!"���ړ�G�8�k+dz�ۉ�Std^x����ïd����c�L[�&L
��{r��^�TQ.	��O�~�&�iֹp��ե䤖����xf��Rku�����Rћ� ����ٓq���`����Y4;��3k;JC�������S>�m�*��N'���0���ʗ��"���&6x8�o�l�@�㹯f�k���nr��؞,���f�2~sÒ��o�İ�?<�!ю ��/7;t��J^��� �[�n�ytY(9~�+���]fA�97�T�ZR�A�6�8�s�������RJ"ӗ�;an�����Xn���������LWl'����9��V��W:�E*������|�<��(�a��T`�}�ْ�|��&&^,~���j.� =z�s5ڍ���PfQ9��/�
��������~���>U�֎G>�6��y�p����ՉR��\��dN{��X�^���I����,Wޤ� �<�����T���MY�VR��4\��A�B苌�)�p72��5+�#��r��VjQ"�Н�γT�cTʸ�x{"��{�h��;(��̜P[��S���HJ����̡��f�ً3t[��5Sgf�~Qj8Cs�/��%��?���.n��p��Z(&t3^?ފ���M�l�<GyH����$�YlΈ�&�K���v:��Y��~�mWyc[�y�1f_GM%��+�T~�7�Ɏ �� �OL:vgg���EJ��L"���^���?+��Q��}Ebh�3̈́*-̄-a�~ʁ��
��/�^\U�U7�*�nK�?c�g��!	H���8N������k�k{�M�=�(I��)?������m���AN�z��K��s�$S�4xZM3�tr��S.
��	`S��{�V�Y*=\���ͽ��;i7K���-�;�,�z�GDU�̖��X��Ab<V�RK<���2�Jw��;�&+dEN�W?�d�^-��ރ.dN�A6"���-o���	��@K/������u�}W��O���4Oĵs���B�?�!k�^��Dp VUQ��b���2%�*n����l��'���*�j� }��U{XLb�7*���&]d�?����]x'�ɨ7P��<�I�,�k��QrK�q�2��)@8n9X���A߹^A����o�򘼐.�cH�jhK���4�o�O�lW9"��y��O�<a�㿥�&zló�ق��D��;�7�yـM^�i��k�p֭h����H��=3��>T"�D��s~^��gUy�C
�T�
Dȁg&��2�r�gu�6E�\�J�Y�eE*�?p02�Y��w�n֑�>�Y	S���r�U����Π:��>�\�d�!�Dڎ���Un��dXe��H~�f��^s��o}ta��o��,.]�['}%441�<$N�qPx��:��Q$.\�\�HJiMC�s���M�ن�eκ��Nt#?t�s8�wD`�g��EF�='V���)��٘��(���Z���Ƹ7jB2P>`�<3�=�Y�{<Ϫ��'�P�R�t�$��>;b�&A�V� ��k+H~R�����&Cͦp��Q ���7�0�$�{V���϶����r'�2�;2� �^���Ȇ��=y�46cw-V2������S4}����
�,W����ϴ� ���G2�
j�YBU~���u'Bf)���GJu#����f��:�ǿ)�1[Y_5���Q����ͷ�����y�p@�@r��\徘�Z%��9-b9G��-�+V3j'�O58W��F����U�k�&��PDH<P��y;Z�\u�n�y|s���˲���^V��~�"Q�9A����QI�)&[�
�:���M�����xqȑ-�� ��N�S0t����`���.E�g�?��I�$L������;d�4c��,g�����1�)sp���d�=N��_�m�r"kXID�����c}X�,���&�0Go�* �Е�$��h�PkFC�u$�W57���D���{��,H��T����:�;,�vg�@��'�j�ܗpcddBl���o��u��b���fŵc�ٜrn��aϜ42��x3Y�b_k�4\˛M+`n��f�_�lj-���O�rd[@?<�:2����m`T�冡�˱����ztt<�3Ml�d�q�v���7ǅ�s�})�3°VK��eH@��{�����ҍ9�\��|�k�@����h:��'%3Ie���cE�� y�ЬYl�+?}���<���:��H���� �3Y|K�4r�����q��"*>R�ٳ���59�Y�њ��M����34����u$�ɦԼ�n����X=�ġ�R˞O��" %�ҭ�l�z���+E�AH���R�P�D�=& ��V��$�s����VE՛9����V�����
 +���-:�p-I��Pp۟>��':	$�C�F^���x�i᧤����X���5���	!P�y�[���#���f�+�H#B?	ػ��/39�~��]%vW�z]>nh8���?�AV���ޛ~x�P�t����pbW2�|��Ǽ��2�_|�#��S�e���~��;젪�������W��c=7�ow=cJIP�tb�n�LL�0JA������!��I�T�כ �>���@�RH���D3�N��Y��a�A�QK�Yw/˗�&^z��.X�4��'׼:�SRE,ƭ�p������R��$��ͺ;nܣ�L�i����U��-^�9q꾕|肥���r�j�M��e���*��Y)o�^�S��3=�}��$�Vzj��$D��4 琞p��w����g�eݩ&�lv�l�����k��K��"lR�̺C�1275YGs&�����3Ot�Tj���1�@�d��k �>��P"~��u�d|�����MG���J/��r��k��n^qZ�a<%�s�k�{Y&�,{���ђ��E��.�j1v^������c����K����FƑ|�1���V~"f6�6���1��tc!V�sۮ	���9����-��Փ0i}lc��鹡ㆼd$-�x��3L (���Z�1�i�}I]�8̟��(L�B��	?��S�k!Ȯd�Κ���>���S�I����w�&�-�Z�� C�נ/�ٲ���B7��wN���V���@��;�c���+�t�;���Ҹ�J�4��)��6W�Z�;l�xan85�p���C����"d�$.t�1{��Q�e�=^v�+IL7 �"���Tn�!��GE@��0s,L�Q��z�8�\;^�؁���������蹗)�t����M��m:�wZ��|���N��V�V�h��P|��;&�ݙ�i����_"��4|4���)%�l�^3k'�`s�Y�Q,����~
�k��ak��U���r9��+�u��8�#�����MuK�
)%-�(����z��Lȼ�ѾM�_�gNi�^�9�rvO�����q/�z22�%b2�ͿRM�.�m1%3�n��T}V*�w����nH\�lF��p��B�RG
tp�U�rސ,�ذRU����EE�����8ku>a~��	3��?3��{I�_��-�UO�[�4^H
8�3��:�bbX��gg$9)�h���'�^�<����_MFh�*pA��Ȼ��p��b<`�]Ǿ����dHD[��O=�)�,���8�7�Pޗf�-�@���+�+���|��F)�r��W��x��z?����+m���h.������Yg�/�W'�`��|��h!ϼ��|� �n�owY4���f
Rτ"��m�7�S$��<���HV��{L1{� V��m���792ŗ���b0��uY�[��aū��x��cV�i��u�����W���m������x�!�~P��1��0"��7Z7n�"�~����P�kj�*HIKgÆ�bZ$�͍=a˗4���厣�Gp|t~=k�����&p�kd���E����;��iB�#�3��|Y�F�w���ƣM��*�ETK��9�I��8�^��Yǹ�)
�66���8e�xy���*3�lk���%����ا�Z������c�}�����@��[&�>�I!T���5����Ȭ�xU�L��;jۄ��ط!�D���CX�zI�����+3�mM����Hw�l��O-�E��o�S�{��^�ez=j��qt�Kw�� �+!�,�H�0$y��<��3�]x9;Y��Ay6D�S�vO�cS��0%��ˣG]Z%��]���_'Ұ���Ԁ ��O�W�H6���gþ(� ����f��9���U�G�/A\{Bo����tց[�T��ܦ�َpV��d�2AU=m։���;���uB�Pi2]� ����%����])HmD=�I���N
�����$�HH�Z����
�g��{����B	��`���{#qO���J���	�䙼�=b�I˭}=ڨ�he@�%��B������݄��9+TF����yE_k���i����5z��E|�K�V����0b��ma��j�BvHHi����6�~~��Z����}7�����k�o��,;�YD�h6�j7\�{� �?�Þs\�[��%hixђ[PdiU*�6l�I\��#I��#�Z�Gy5Y�����x.�ǲ5Ƥ�1��o�U���!���c�x��z?c��%D�$�@��r6�X�" ZU>Q�#�WÍϮ� iH~�V��y����P���0���6��Pͻ��2q<����u��@��q�I�=��\{J��������	���ڽ$r#��H[	�훽��eR���ޣ1�x����I<j�R�C�#y	]:�h�$�<z�t.n�,W>��!�p��}�L�H������!�)�|9v�9_�� ����x�=dIP����G��wC/[�<�%v#�J%�37X�)�I}�^��<�~�$a�S��6�D}�G�Qh�8���� �B��[��ao��U��!RHLOt_tbBB��һ�m���E��^�k�Q_	-vb�;W�7���p�Ss��0���N�Z	�n��+j�����{����P��Ȏ֐���
�0O�<!t(�Jg�X�^�
"����-nT$�V�MM����TS��
 �����zu�x�(���]���V��_��*�»�_�T%�K�ߪ�P����J��a��ǆI�S���177w����uw��
%�����M����J�<���F�H�C6ԝ���<���`)ԍ�ge��Y����1�:Z��:�V�"|�3g�������7�Zd��B�|;R=e88��$��O�������x��Ȕ�({��J�X��0���qZfHc7/���	z�H���Z[`E/	]����`OQc��3�rـM�j�gL���ţxG@줻_"�z�q�j�tr�V�u|�)B������~f��-}��N��_+v.w��F��:���k��HJ\!bU�A������n�q>+�����c��-���l�����!6㥪\�8j�"Z"��UA��R@���g�	�0��Y]-�Zm�2q�����t�ڋc2��/��먠��U'X�W�����X�g�?!}�(����(�&�z��1>��/���{�@0:*$\�[�_|}Ҝ���5G��@J I��6���fЀ�����5�>�:Eg[ɖ{���%��g��jZ]���2�9�k�N�2����$�"!���8c��e`�Ie��H}i|q�]��<��v��X��7�O�qOXD���F��US�GGJ�n�-2�4�x$$�}V��y׳C�~r~l��G
0ڠ�ѡ"`�)U���1׫AV��%%j���H.N?�ڒQO�t�yź=���T,:2��+�H�ʾ�����8*����X(�6����v��j�1B3�^'��)�U���!b�/�)����r���j�$�)Z�yWQ�H��N��7���^9��P=p��8�i�JTΜIz�K%�A����ڬ7�5$Y�?^J�Žr��y���q��ix�k���A�"�0�o��+�L�A��,Vd+ly����_�����M�(c�ￌ�>�d�fi-5k2=�����9ܧm���qӳP(	8�@�m��gRP��I���e���YhLQv_�+k"�γm�X�YZLA�k0�1�&pp�:���(*��1�$��l��j?g����	@����BF=c����^٪yB�G��Uxq�;Co��3B�㯧�]��5��Y*��ʡsNc�f���b񲑳d�#������MZ��I��Ŭ:0�cj+���S������p��k�<g���7�|Ul(�v��r��7�Cs�F��糠�n�}�Y���(��}e�X">���Y���F���YW���}�X�����)t7��|������	�Ne�rd���� ���b&;۸@�L&x�]oZ|��A�\]V6�1��46�D�e�n�����dϠ��I_�,��[�ôw������:�ޅi�FZ@��K鐖)��$$�$���閎���!������^�����kÂ����~���>? d���6-.��P��g�	��x�k+�p���
k�S�]�p�N�U�&��K�I��f��S5���;����"�խ:1+���eI{;<���/W�@l��1Q����Q���S����w���^bGSI�"_ż�����elX��vc�g����8%���1GS+�Զ;����j-�z��b������hJ
�
W�5��K����}	�����EU�=���X}�L��8����R�
��U��e�ɯ��
!�s��nZ�Ƿ����u�F�}J�<���U���\F�v:W<z�ʧB�:/`gW���wmi��f��WW�a=��|3�����]�_XK<���t��p��]d�:���}n!ӽv2�3��Ba�ò�PX�,����zj�=�̡���2L�R�i�)6�����'�\Z����4�w���/֨���~=��m��BC�&�&��ܚ�Ȧ��i0w���Lg�{�:��8�(���tΘ��Q<,)8��̽4���NF�l]�<J]9���I���+�ɥ��������%���1�6�����݊ؤYe�%�CGqOm��g��iFZ�6�K� X����M�O�%�)��g���"�����n,RWp�_�2��t�h��5�&4;$zܿ�W���2�m��	+��f4pܷ������(�p���]܌�5���L<S-�m[qV�Q����V�2�S���h�?Ľ��S�c���"U1Cޢ��֕滖�:k���ũ�$��Bؠ���x3RQ�R";bۉ�X��#����_R�2����B�bJt5�������qcjoE���z���f}_ېښ��F�
��f��N=��m&�z�0&m}�ai��(�I��ͮ�{�/r�2�������	T�Ʊ����\T��U5c^��w[�����ʌ��5�Z�w��}����.dP ��O�f=���0��:If@��pO_��7�7<��)#��5�ƹ�w���djY>%�F��;>^쿒J��m���iɩ�^�ݴ�;=����������J@��D�16lo����:�E��p8���������^��;������)se>�/����
1�0�5Ql&��v }
�<5�i�f=�v�ݬ�>Ϻ��)j�W"���+_����gm�§�n��6 ��>5;u��E�4��g�rgx�6�j9K�l\YFI�}H��p�f⸾�1f�:�w<�۰\�����q>�����������+����O�;��!�b��d<�_i��s�+�9����0�豠�%,�C!��]F�F�Y��-8�}��o���|Ν�>@/�L���ŀ����Q9� ����,N�5}�꼮Z�`W���.�Ko^�ś]�z�~Z��}Q�`���|Gr�x?K���m�J�\(��20a�O���|}d���o:Q����ҹ��c!3�p*�'���)��t�w9�ߧ�50i�^�m��3�H� �_��
�O�LM�1��:��g.Q@�v�p���U�li�n�%�����S���x�7��L�1e�ֱ�ZB��������":s@�5��I~#�Y���f�N.��bO0[6�z|����}���R``۫1M�&qnC��~���U����E8�2�,-_�܁g�|�O�mF�~�r(�K�	��"݅<�̼�V�F�b���̈�������f%��l�J ��*���m�W��z�rC}��X�/��0Fv&z��U���#��݃����+�?"������+q;��&���A���nX��Ĳ�h�x��l&F�|�D�^|j�\�S��C�y�����e,��b<�T v%)�,%��s���-J�Y����_c_t��b1�Xk����0�	���p�*"��%�������2*)v������#���m6��o̭�nG̊)(`H�j-"�|a�����f,�|��V��ETP�xK=F����~6�*g|$������A�F�����#i���IC&f��7�^��9�=�-p'5e2M�J�/���$�AǧkM��]��&�L7�lH�N���s=�v��g:c�R������qD��!blV~�vJ{_J�Lj�S���C�7��2l�=�5>p��xm�̔���7#�����@|��������;�rэq_{�_������uD�J;���[���v���k�e_���	m[�=ᬐp�%�����eD
�e��kw�f�uPV��`�G1��LP��>a�/�y^���Ƹݥn��|���&�M��֋��4�?��~+~���.�����#�ZuHsp���um9����#��/�vI�P�К��<��RH\\-�_�����؞�W��5{0w<��yH��U�jT؜HL�ʏZb%���� Ri����'���Y��mkT��`��(�&U�|�f�7��1��dxd�6���]��J�8mAfB(���N=�?A��5�-�����<����zE�P��Z�\œ_�@�_}7�z�g��+��+�[Sz58����V[��BժRPo
�<u�45[�G4�7Xk�S��c�}	 ��Q}<>����������u���=���6SլűM�ݮ~��犕ЁUG�b+jB�Is�p6�
��X�cKyg�L-B�Xgzϣ�xH�W�����.�;)���2B��G����\^Wե��C�%>���kc���w���F�yKnh�>dg��ٙ��=��߫�C��P��ׯEkR+��;�  �S����M*׮4�Q+�C�{�袜�6i!�sy�W�u{j��X,Y\-@7[���6��iK~s���+󖫵�6�-����'�UȘ��vl�ؒ��?#�/�;�"�~w��ؾy){�Ir�Z�!��4C�{���қ%��~�@@'�a�s����o^RL�\���=�op�����&�;kT�u�w�4��`�c]b�yOOhg�B���vTW���4r5�_!�Hw��ڒ���6����A0���[�^A
��.kK��ұ{�0�:$�V&�ag�����2��kt�po'���gUr���9�w^#p��p�i��R뻳;�Td�D�9�F�c�(��Q<�*m:@����c[pj?o�ro��b3��/���5$J�V�����n��N]�9�E�/�o4���ԐV,��l���U^��kꞻmʭ5��إ�,��1=Z�`X�v((Ѯ��hQ�fU�k��A��s��SPh����O(�{�,��F#���Fy��c��j�����g-e#vK��k���	r�#_/1�c��õ�1�y>�|�(�P����S��I��6�O�T��1>L�#���6�S�{��3��J�V2��f[p�����᫟���j����tFg(�m�/�ˮ����Uu���ގ��2���E�n.��+�DEۯpP��_<�ZbxE��7k_�RJuo�՘X �'��UW?7$BMzpMB�[�rT�fk����������^<�hJ�rY�d�!�q`����a�4hd�I�U�m0��D�@ϫ�-�	y��m�|(�㶔�����0��m-7��u��:NQ �8����FX�lrk�����193�{�V4�|��zS]�w�1!�.������Z@9�
]	�j�A��IQEO�b 秼��|w�^J��@��N��0�"��wv�/���W�`ln��JV9z�ZJ�\��,Y��?�W���#��uR�e�1޵W�:EhQ;EG���~��K��;��
۩�E� �����~)uگ?/�� �;-:�&x)L#���X��?���jr��B���ݹ\��!�s�a%���;xxs�D^��感ԇ�m^��|���ccޔd�4<�61G��v}T�F�u��Xz�
�a?�̑�U[�x�AQD��3l�1I�����	!Y���:]��߀��_K��Z�$�mxjb|nM�7���&፥��k#Čd������"��Z�>���o��4�1Zk��5�ЄN�ۮ�Qv�2!LF�8�C,^*&��W<�5��,�_�f�����ӂ���I6A����Q\_�Vۋ�$!=^�d����1pTo����/u����
_j��.t$�%��zv࣋��|+����X^Y~��2���W*)c7f�Z�c%�F����i�:��;u�1L���oJ�Rf�VJ���^	��wx�6T2&:���|�0xh*xj�u���A�3��@�S�b��f����;�>�0E���uU�Y����!<��W�����)��~X��p	�<4|1�Nݎq���@i��؊4����k����`�s���ZL���6K~���m�.����0�/Eы�F�DJ��; LM��P��=��-�H&��JCJ��o��?���^����aK��QFڼ����[Ip��!��/L����]�wo\qY���^��:zg̰�X�$mmͬ�SK(7p Ӽn
���|���l�o�G	��*qj�<"PK�Z ��T���"��%ʒ΀���9�#a�����8�#�ah[�T�I���=�6,����Ypo��-G/:�+�d������-�Z�hmrɺ/P��^����y���T_��{��N@:�l!�R�����mP/Y���vV	���������@1+5�����uw3$x9S� ���dFF���;�;����lK8x�.3No�Bba<�ϒ�~��������7���E}��;8���y8��{a�.#�K�6�!��}���qń��<�
'�8��%�)����_��ب:]Kp ��oO9����4��&]p��"��A����dv���U�Ҧio�|7^����N�2�
L��݂Rj���?A���Mh���o<��)�ߊᣮ~!�Z���j�]���0N��S��B����j�~��a�;?��[G�/�7��O�Ku�Ih�LT�z� Q�Իc�G�T��{O��J\=L�UP�@�/�f�98�;0��"&��s�����́#�zi�4dһ�N����UhQ���H�~�G�����s\K��
���X�A�.��n�����5�'���ݑv0`^���Կ��(~3�W!h�,���e]�o��8�����Ҭ��ɆJ�1�@@��/���s�c�m��)�7)�OP��toZ採���86�#�UM��/��X��\봚�v�����hH�x��3�ʺ�����^N���GA�w���h=���2���?�$bP �7/+��<�!&���}d��VJ;��'�c���m�F�П*�:+�~n��/@�m9&U���l����H<��Hɲ�o��*��,\?ۂ�����/4^Hu�ĚK�4P�C�3t��C�6z��vVQ����Tb͢��N-��"B�8~��;ܵ�IxL���G�|�C��<��P��ӣ���o%h�/�zD�9�
(��붆'g'3��!�b�?mp��J�ٳ_1��h�3���S��d��%{p�����8f��k��=-�NW0]Wk��b�|�� �{�����\���F�2X:��/s��N m�4b��b\�����h�;m2:��t=*����NM��|z3wZj�������[�ɢ����̹�r����p���h�}�Ϗ��,�g�J�F�'�:�5ml�Q��M���F�4,��#`lX�5�e8�bN3��ᾪ�W��y�:��YW@���*ke�N�|�@�?w$�OiP�SY5�z�H˔�-\č2��6�Z����x���`1?���Fo}*���ֱm3�݈7;��j�0�Ҳ⯷���d�nY>1�J�y��s�8C�'q�ao,�w�6����1^<{��m!��œy_���aYA��Z���
Gkv���+��8p�����C�:Zn_8���~������ �>vd�=<��!2��`�D��ɸs�����߉�5y���?�©���tkЕ�һ���w4A�2��m�m�٨�b�6��
�f�5�b�����Ryk`����J�M�?�拞���`)+B0�h���b p;B�©�����}t�n'�ylkql�(��-PqX�l�m�K���9hsR����/�.��|��	�!o���@�};)T����S[�>fJXlN4tګs3�T��Ϊ�s8"�UDBZ��kj�ß��@��ϛ�ѡ98��Y�R���`bКȹsP���q�6Ӎ�D��G�J?O�#��)+xa׌�@�����ep\�9{��&1Z�������V�gL�2'�rL2I��TRQ���xo��.��F��&�uM�6o��w�#5�E�lJe\q��,�����i�<35 �F{�/%���ծ÷@p�/vj��nf/�C�LO��	 ��Y�/큈pf��L&�+Tu���`�Wzk��ί�vO߃#��/z�f�I�Y��٣����>a5�SO՟KLN�>��=�%B��d��'\nP�c�Eb��n�kT�9� 0�n����h��x����<�\+�(������g]tBc����S���t�K��}S�ˁOq ʴf��>n�1v�9�蒳�TjW%�y}���*-�zFS��g�؍N/��o�㰮�(½�:�<i�9��������y���e�`6��v��x%uʓ��G#�2� �/�jf�Q��T�#.�a.�\2E��f��U����б�A��Jl����eL[bIL;r讲��p��\�-I0uXz��A0z�������ë�l��kF����<��^�=�,yf$�{PO�U�Έ��O֑���i��?,	:�b1��R�U���n��{� .�uG�|�Z>�\XJR�!A��=�dh�tG⹙K<O ������Z���Y�v�`,���c�rY����BQ�&L��2�:��{��1as�/�ݔ��F�Цn�Mj^$L���=���͍<M�@Z�3O@��&Q�Y�����r��^W�q?�������B�2�O(�������p���ɺp�	3KM���y�5�����e-1v1���Mc�,�y� �B����9�jIJ���mt��u
��f�_Z9�[m�Ʀ�Q���ו� ~�ٵ�t�n��g?���	�P���e�Y0!S�J�X-�ڨ�����dg�M�Z�==F���B��e�sI�ҵ�������vq��⍕v�g\+�H�N��ɻ�^4g׆W��R����ۊ��uX�2"���٘�k���=����2�,��F���?�*�ڰ���Ϯ�O��{��[iП���v��[e���-�CA�|��}��&`�"İ�B@>�$��[�V��KM�i�ȁ�����6������'6�q�'�B�kA��l��;��*'#�b�xţ[��[�#�r_�����3�,�+��I�i�гp�y^D�F���{J�l:
���[;���������z�D��y`�
�w�Mv��;����U�V~x(�?�Z��^�������Ϸ�^���ֳV�BFg��O��p�*�����s��Z���r�+��w�30x��Y`��4�¶��H�,�����&1��c�����q`�"$��#��fZ9W�t��z��&��i��ÁS?��fǵ�S�8����_-�{o��@�[�k��oh0�{�ݜ�n&`xPK��1���xei��elJ�X)�|�e��'Ã�؆>w������2��v�s>�;-�tީ-UgT��b�9H�ܱ⩉���+_G�Rm��mJ2,��jz���#[,�4���3K��N��bJ)پԶ��	Lh6Pc:�I/��n����J�53��S��k�?��gСg����ڊ�k�ދa��'�ߌQJǶ�n��=�v@ ��#Y�U9x�~Ӯأ��RA��iSR���M��	���1Ë���b�4kߐ��^)l`��-�	C/�P�-��\r�Шr�$R��o�GEb ��F-�Ջ�a	���Hy���WK7���R�R:L.���h�-[d�^J���N�&��y}���D)^Aѐe*ܵ�*�J�6������J���*G�/��Ƿ���d���z)(���Ѕ'�S��ț����E��g�5	���;<<�g����U�����m\�1�FǦ�.]���R�k���*�l{i���s�>�5��(��fy�T<��^�a�E�g���1��rZ�{�
\�B�L>h�X�B�$�2gp��SGo�ޝ�n�s�@��5g�ԟ�+��w$�`�O���:)
�g|�t��N2�ʵ�ﰟ��[���w'��͆�cJBR�%m���o&�{�u��?���\�v��|��:H�l�F]k��vF������/�m��x�H^=n	 kݓ��ѽ4�k8z20��*�.�a%/U���┣yw%�����?p��������0�����Tm�wwi�����R>�Sj����O���۪�aԐ�5eޝ�o&N톽F4�U1�1�����	�H���Ǜ���wH�*�:���zo/�%���o�FZ�$������%d]�/��_e��;�;k�zg�aU�18�K���7�޾R��V��K�B�qj������Ahv?P.�i�����n`��v&v� �^�����}9=��a<h
�<��S=�>W���[ d�[�t��n�{D�Ǯ�&�Ӄu�M����>�L����%J�V"�Vv�.�T�d_�ʒ�J�BɫOO^��L鞢�,L����?wn�@��Q��?*-�	Q���a2���s��7F�in&f'g.�35UÙ?��lE��^�rTMP������i:�!!/Лf4�N��8}S���rHp�L�픔�W��<��ܼ���uG�0۹{Y6w�_���ޗO�������)��V�}�,E���� ���I����硧 ��ىv��Q?�A9d����=!:�+��� RP���y����c�&�0:6�I]���C�^��v�ʥ��{ҷCZ��:�@&�R�wr��'3}�P�i��P)��gh�� w�jw%��B�����M;2%�{~J����װ��*k���o��)��F9��&�FF.���P�+G�!���W�*9ܹ[bG�|�a���C�0�䮿�	������OZ��F  E���ؠ�{�c1��'޿�(�LV���O����` ��Q|�(�������ehI�!z�N�W`c>_����ar�?Y��W���b�(!7�0|#Z����+��C褷gMk����v����x��W��!ӬQZ$K��2���ԙa���zcR1�R���=/~Q���mg�օ��{���\!i�(��U��𯏙��h��n��ES��5i|l	X9�k���Ki�L܉*�0��ȹ�D�iŨ|�6�������S�zٗQc�4@ɱ�̹�A��2c����0?�/�!�*g���5t=�9��ܓ����̔4�ˣF�hN�Q�7$��k��v��vL�Ȳ8�-
R�r_���xFU����`廽/OT�)��󥦁A�ǖ����:���gL�M�&��I�0}����G�ui�P��`kÑ�3� ���U ־�k����e9�/������y�����=�*�R��|r��V��~�~9T$�����3�����;�0qA�j[ߵ]ur�M�fl�]�5������Cٷ�y��?�/=�	V$���%?��7 �:�̜'T���~,�ڵn9�GȾ�V�Ϭ';�����e9���&���# �=�sf��a�ftɆEBb�>�=t_�1ci&�B�6�
#�\Ú���B@v��"�Q%/�H6��־'�Ɏj��N9J���v��|G�� '�6p>o�!!���޷���\勧�(���L�G?��y�"n��RC�GV�N��n_�ܔ�x��P��OG���>D���Q�,�G�S�*)�/�=��y'Y��Q����B���� s~Un��཮���H� �_.)��9�1%��ڲx�,`yO2=�¥����K\gMD�k�(⅏�Ԟ�V��P���Y�;���r�T������S����!��f���it�b)���v��8���P��iV�+@/r`���¹OJb!��G{yT��+�?[��i+n�m|��l�i�z�4��q��[/
��c��;H���E��%�[|�γ"�����YU�5���	P&a/$d@�������0�6�0�xj?�/��8���G���*_��kEiMԒ3�vp��	�����p4�j�В���YXb��|}K�l�ԝ���@;M�����j��b�p�n'K��	��ߜ�y�Ɗ�-�{����~!؀SX������'����(؛I��-�W��;�'5��ڨ{���Z��[Vp�h*�<b~YW�����3h�f"�1��S�I�.�W�+eKgX��πo?.�HM
�d�����4Jy=�$���r�y}�/%�!�g�u��߲��oZ0�d2���3>���^��4
���O���/�ӥL3��vV��������Q�Z��٘�u��x��7�#/|Y�l�*���yyB�i�~x((��p��Opdds��Tڽ(��k!��I��RO� 4�B=�ΙZ8d�q����p�*�'0{�2@R��ՠ������km1�!e���[��<���}�;x���'͖k���0�6[ZuI 9<MrP^��B>�c���C��Y�@W�/=����P��2�WR�J;�ʀ���j{�e��<K�x'������rh>8�r �ɡ��$	�����������
m�Fh���K4�9���#��Bn��]R)���p�*X�bMv�.�Cw����#S���cs�gG��m��-�=ӛG �>�E 0E�=y�5=���a�ʦ�3��/�����k��Ji2�R��Z{��dM��c��u���	껭�MN��J�8�%�"�&��v]��&��Fie�[�f�_��k|�R
���p� �#D��R��&!1�� j����d�V������F�@������z��ڥ��m�)���67��ߵ/��;),V "��p#��Չ�@��zQbJ	���Iw��U������|�����l�S�9ܘ���o=�L쬴�C�l��W�����	�$���<|kh�9���@�Ep�Ĭ�L�~޸)@r�����S�t�ќI���S�W��Tx�"d
G9�����1[;�J=���@a�<�����r
1���5ĭ�7Z��q�Vom��tn�4���w^2~���X��;��)��΋ٿ�	�M��:�'�\6,��՚/KX�8��C���v:����'v䩷�c��H	d�j��+$Zğ+���g&����<��$�L���~e	N�	 �Ψ�Ȼ�$����ގf�1l�q�A[U����3y0��p�֘[��84+�ZmD�.�?J����"�#�+�-�@�&-��G�0�����uθ6��&����ڑ��C�-��ţ���Qc���TXi��WR�_���G�w���&4�8N?w|i;�)y<^���u��Ħ��䚖Pk��S��L���X\o.Zk����<NJ����ֶw�dN̝� q�-=��q�XHG9O8�J� Z��l��y�۝/@V-���桞\��7�q�n����̷Y��qk>Y�L��6�O./�2�����h~��pX�=��E��wxt��o�"b狨�D�B�U�ފO+[m5)���Q뢼o��U@P(&h-��$ξnPK\�` �.P��>i*��W��ӂ#x	���NC��^km�8�R����,�
(�$
vIP�5\ 8�?�������`��Uۺ�4�ib�?�˸�$���OJ�xq`Sz?�o������%++*>��)&C�M��7�R�r�v����8~��~�<��}F�0`GR[�G�kPK���e@8ֆ����H �bqrk���P6�ϓ��0'��3T3�^~�/��`�A�B�ul��d/�"�E���k8�
���幩9���5�޼�����gJd�Z����xxM�0�3'���*"�������0^����x�tn��sJ~��&;�0����Z�J�ۢ���i���)]yE�ua\�zN;����\\�{kr7��Q��E�0��ݴ����	�n3R���l�S\\�um)�/��N����X�Vj[�Nv3R�A��e�d0A�
�d�إIo��^C�u��_k_M�����UYTM��wX]�q�O���y^2���P�I���w�2�B������ݷh�S�NP��LФ��-�,[yɊT ��+��l�ڪ�?��2>d���t����Q/�!���E�Q��	\��Uq-��E�K����	��#�C���m�G���ш�^��e������F���>�����v�7��#���;:���j|}\N��ݟ��Y��1�����v�Ζ��]%v�M����OA����*_���,Wc�Wo:�)&@�N\����_\�Z\p�|�i���駯���{�4���R����~{7p��lK�P�O(Sr4"����z���)j�v��1�J���oom��޷�=��� NO͛�[|�M��M���:�˜d�lpB��;�������Qh[
{�l4�����Ǫu��?lҸ���,��Ƣ��vL���Fa~s��!�ZU���Y��:XΏ��{�A�+���&ﶙ;e3�]�}��}_p]�l��O��f�א�g9s{��4�1�&�~�Xz����7c��c_�K��r|o�ƌ��@�`ٔ�����L�<��v���3�J�ͮ��� JA�w�о1#�)ݗ'+��2&�N�mb}�W����k�q_�V��g�t$�N�[/5:OؓZLH_J�R��A�f���j��&�{��Q�$T���͖���'uH��/�b{���؟GO�U~�x�s^��!2E��Go�G|e��S><�&�*F���G[�y���v:dIg:��1��Ý��+��T��/�0�����Zbh��k�C���Y[-f�q����B����Q����3"L�J�C�X)t-�A��lO6�`q"(#�Lm�ku�����V�ё8U*8?_&x��^�S��l��WB��.N��I 98�xw�g(l-�c`e��O�t�ْ�j$�ݜ�ħ�L��/����__�g���H���O#%�Ho���}��P$�u�:�A.��P�Qe'4�����zf=���M ��g����Y�@n�M���b��
���M� ����(V�,�mԛ��8ϧ�-6����V���b�����N�d����5m,E]3��{9���a�CHH���s]y���a�B���e:Y���pfP|��Q1Ǒ�`
*���������WD���#���V��xV	��m�ᤔ���<�v%�h��Y���p�.�[�0����_��`ҋ���A�%����b�1c�x��]���qZJ!�Po�[(D5����=�!E��׭����%�sׄ*X>Wny|º���}�&P����7S�)n�0X��)�B[@p�W��I�#zM�\S2v���5��Ul���W�;���7=�� �&���(qj?�+�vT���?#��
��YW��"��ӂˈ��~b���ԝ�IC�J�}��Vv��r��	�̀'�H!9��C[�w֜�S�@�<1�ĘO-������̂~���)���S8G���m%sW��x13�.A��ͥ`�;s/�Gq���3����g��E��U�.P��m��_mB��V�=����c�f1`�YPY%���]����2�>��
^�WI
��[i�����(2�@�N ��>��7bV��ӷ��C�����{K�W���23�����зl�-���(E�C���?<���J������b�*3�͑��,����η�q1�j���@�����-7�|���,�*� �Zuΰ�ѧh����:;;yw��sh�$���r����a�s����?�@�%��4Q��Gg7��ߜ���L����u�:�v�&�����.^������=r�;��q?>�&�_���.nY�"haMۑ��	5�tP��	6���������>�/Y�c�V�^���6�'Gb.����1���AӤ7^'í̶1�N��i-�FeU����X�&�b)U�Y] �l�?a�+���W��r���,ad�CQň|���"�q���� �!���K�U����@��"�H��m���E��s�o�m'���_�� �j�x���4�\�7���;=�[�������Aq�b�N�������4"��"<�����C���O��@L
?j���9\�;a���+���!��aJ���Nrꞽ��OF�eZ�h�;�Ż	~A��{
�^1q�n��W�9�s��콕��#8��:>5�fy����7_HL�Lx����l�]r��m��XkCY:���@�5QtgZ���f�kDxb@�uR������c��*�%��N!+�JЋ}	,wQ� �E��f�ԉ��tl>&1ͭ���$��k[��܅`����C1Y�\6�����;�c?f�h��T�%�D�N}�!��_e|�sMY�βlZ�Iyt���BQ1Э�������X=��p�K����"�I6o3������yJf$�xļ�Q}����x
q̔0�@��ԑPM�m�'�y���+�:�GY�A��!�W�Z���\<y��~��t��D����t%�,~J���I��c�`��Fuq��H氍4Q �i��'�{1\�K�r����� _��'~oϛ`3�᭝+o�KΦ�%-Rp��$�����i��^V��┮y`Ȕ��@���M=��A��F����R�� 2��6�$1���ըi65ER�i���*h�:A�?��ڤya����.���L��/7�D��[����L�@0TX[��t
\˲1����*_��Z��K���^ҕ~a��M�i	�ܹ����z�9˸�z���m>1�x��)�W����ЀE��و;����Y܄Ѳ�}�3I�wy,w�({��{9�$�r���$��o�E���s�kEJJ᭮�\�?��5���!s��"];�l�۷�"yQ����C�i�O���V�ޜ�X4����I�M�Er���1���Ҕ��������s�&�2�b��ο-3��������	��-���A�����C��r~~���p
%��]2�ĥ�>a���%+[�{�pu'��4�	��x��?	��5�_�Զ�KQW�Q7�m�30���i+�;j&Q+��=�H5��rs�x��0�C�z��0�v�$r��W��s���yL&��s�������κ\X���7^t��/�kk;�[�z$b�:�t�[\���o.�	L(07�=ފy�bqj�� x?@&����4�F��ȩnҮ��w-��*!�:�,8�I��UC,��y�?�w?����r��:m�Es{��WCv��t{w�c#�Y�<���l��s��߶�S�A�<ռ�x�t}�Au�X����_��<�Q�3����/p�t�\�%M~�^��"U>҇zQaKE�����s�xSv!�{3�7"���`���������$��3p�zD�g�"���IS"q̱k��4�!Zz�5@��khG�!�L�u̈�-�m��� ��-�,�����"�RP����Q6˨���$w;p.����Y[5�r
�Yޠ�B��.��},Y����}�bh�&��A[[����^-[j�x\�l��eܡ��vlT��$��ʖ�J��J�_2LeA�ek�����R�=|O�-&O~���q�@>�a/������*��1�*B�lu�Qy�6�/��:�ɕ�BK�S�dzF?}��Μ>�M�Qî�Z��V&�ҍ��V��c�h*�_3��>ˮ!�Q5�c7���;}4 +(b��L1o��3CHD�9Β9�4����wpz8]<��U�Z�� ��^w�1�Z�X���T_|�쮳�ou #6A�␠S�{F+�KF��/:?�B���l�J�AF�����Y.�q���m$w��C�bC(�7h3��U�O_��"���f���B�5�/���x=�r���hYᇛUl0ԉ=`Jf���u�`V�B>Pt^�zC���P�N�y��Y��M���<�,�]���CV���_�g���.�x�@�`y�����z$[?Zn?�xq}��w���s8�%��������/���m=I����x*���ҧ\�WI3�O�^X��@ ��ST��>��[�w]��E�����3�7��ĝD�����̴W[s>�9�9h�x�� k�;�����=e��B_��'��Z�g���х��o*^�l��x��r#\�칣l���ES���(�x�βyJJ����j��s�@` #�T_���lw9���D��A���DQ5��������?q>��*��2�Y�SwQv�.���%?�~N�\���x���x�3<wl�����&Y��X����=n������Ł���h�
�_C2��U�9.mE�2�T3CI�ێ�-qs��Ƨ��?�d�q���t�z�t���(�7G��u�HJ
n�)��~򲵿=�I������uM���དྷ7o�`�+�G0����hnS��fg�N%<	�q�áO)�L��<��`f�OVB+�p%/���ˀ����9�&�Zʆ�
�(Tbh���-�%Uk�_KFG<�s��Ё4�IG�h�] tڧ���A�����K��,B���l�Xl�j�=/Zȗ\O� �8P�wl�$�}!���Jy�����,e�ep�'9^���;f_��~|��d�0ۿ�ǟP��;�2�iɏ^��p��/ݠ�s�m�Y�]ݴ�ƒ���J�[��l�Ϡnp̝P�)�1k�4>��^ڏ�
ep���W>B(v���z*+ZȑbPDdz��s�}U[�pR�0����c��i��=<�T��,:*��}r��K�Z3�Ax�A��4lF�0;4� �я������_������ۿ;槸��{������/۱	y��]R�T��_��^�J_\"����뭣�~��qP�n�I�[�A���ҭR�C�i]������=�7޿���|>��칟�����g��A��#[�/u�l񖿢a�<ނ���������������J�n������2ݍrv���k�(�4A���ۜ�w9����[N��R�dp�'6�c��/�D'i�?���o����;d�\Q�R8��7J���g�C��G����զ���E����V6nB�� )zoD�nƵ�r9J�h[�¹n���a,U���gG��=�y>�vّ66�<ƿ?�i��_�&�wdBNP�k������`��󋙑����HG�I1��3�T��Mz�$~<�7�f��F
��ŧ���B��"[&7���:&��OgYH3������k�`�Yn<]�e2�֧x�a�y|��+�kg��U�iey��s|���'�A���3�6<��]�8������%IeU�*�1���I���I��"��{���K��F�݀s����36�h^��
�rS��	Q0 ���IKx�s'��_?���Ў���-���<���G6����l��<��{ qa��c��K�F��K�y	7�s�D?TQ˥;"��ׅ�i�]�ӫ�U�k]��������0�Aq+
���擙��O���#������l3[�)EN�G��!Q_<���\8ze��J/>�GR.X�-�{+� |P����U���4�y���R�]���S��R�yͽ��	�C���X'|^>���A(d����m��ǥ��rt��'LqC�������LwF�*3-�}q�n�r�Cs��V��/N5�
�J�v0t���]��>�T0X8��j{����աF�9Rjq����F�{�ڀ���Df��:-e.���%�ɑX�.�X�n�ت�=��\�k�{�U? �Hd<$�7,z5|z-$��|������)	��;;�	��=?]�!p-��ć�ۂe:^��y�O�G�&��֖fo3�w�(�A��'�V�j�Q�1w��� ӆR���c� �Y ���fuW���rI����C%�ԗ�x�1��v���_A���r)��}��{��C5)}�0�MG3�K�E����CiB���
��,K��{����Rf�:��B��v��}�#	���AC���U����K�{��6O�;�V���8��Y� �B{�Kg /�ˡ�YA�yv��d�rb����j�����C�@����+���8�[GM����*���ww����B?����Y˪e����í�Tc���m��0��#�S}�������3����8?� ��Y2��Lp"t�Qa�8ӊG9��U-;$���VlCV���;�Yc��"�PK�ܖERg�
;:"�+��ܻcJ��U�������n��*��ӆ����a����x���_BH?_#+i��&y��
m7�F&��������8owV_���]�s���h�zd9�c9P�#�M��̽_:/p?o����	ؗ7���Գ����Q���`����,l֍s(W4�^�;�`�'������O�/��ȋ�*{���3��*ݭ������31F5{up�1�|��ͳe.e�d�	M�K�z��Ii\YW'*zם�I�n�]�ɣ��Ěw��n�B�1��Uv��+�?�����>}Jul�z�W繞\�vk�UK�)R�/�g,� ƫ=4��Q��[��?��_fZ[���]�|��%��۳��v�ݟ1��/Ց8�����b_nb��~CD��ɤb���F�a��q ���@�y�I<څB�q��?]o@'&��!�-?��'��i����_0���y����"FI�̶�a�k��߂>h<���MTf����%4cZpL�la ��~����6��>�b�RWWϣ�K��gΩ��*����^?���Xx��?�e[#���ǱF�"�x(�=�������˾��K9����޿��AT>�i|W��A�$v��F���,>W����p��O��?�5���(5L>E!ZQJ]����U*��@��¡n5�.�4�����TY~7N�f�a����=,&�`f;P��84���hky�p�H�ÝX����,��HU���3��ڗ`�KA*f�gz��!U�`55���䴍���ư�	,bH��+]����������Kq��)3�?h�yp|~�D�e�M����ft�
��l������M��E�R���4ÿ&��Hg�q�־
�D�[��y[O���e�n)�T�x�w�-��	�,���1����d��N�C�o���R~V�x����9��	���,��u^����+�am�P���[��R���H��S�N�g`ʛ�;~��<L}�v��dm�O��
q�kO{��=h�uf��+7��7s���O�wָZR�0cf�R.�;,�E�j/�f�s�3sYn>>sAG1[6��ސA�o�H*D�rh�J����WUg�����b���h$�O�T�V��gㄳϜkV o�j�+1Xc��z�~X�-���گ��Z�]�lG��<�8Im�����&�y��!���0$�Vh�����6H�޹��K1U��L`���T�n��+�6��(��U,��]y��I�wq�\XT$#��{G�Ր����P�K�b��M㓖z<ܦ��7�Xo2�ƈ�;����7��(�@G���n����F��&�����ͣ�;��օ4����P��r�-F�gn`E���8���U�WH�A��j)�h��qh��N��\��]��3���89r�O�G�f����ru��V�7oh"-�>x�t&�9�p<@uX�_�_���?tIm��{R~M���?g�!׵=
�,\�oz��U����w�����?$Ы120�u���Ih����]��O��@�q�NJ�CxcT�9������G`(`�+*653��8�Y�&o`)M+�
l�>������ֵ$��D�Q~��Z��d��ĉ韶f~X�V��Sǖ��Ȧ�5�q�lq�P�P����%v����H�w�+
L����K_�+v+0���d����Y���T�d��~���I;�\������u�8:.Dt�K���+�^�u]�g�F�o���� ��|����xu������`c�M���{�T),ɪO�������/F�V���j*��<F=���<��?�Jbό�y���ά]��ak٩m)�/���ջ�b��#���
Lq9�CC*�$V�|v��Y�MIf��[ap��Ds�9yΎ��N�F���ݳo�u|���w�v��]_w	P��7�l���Ji��S�31������w%n�q���GT�����)����J3]Q����gp��k�z:����wn)�9Қ����dr`�/+}#� ������y��ow�H��r��Px�)�����M_�3��
�;T�����R�i���t����b4�Tpm��wT��1��f��,�3���f�'�a]e�c��Fm5;�?�p�=�<�ݍ�����*�k�=(;ﾹ?���1�!b������j6�S��f�f�E2�k%c�[;��7]8�f�z��v��r������xg+[ �`���,���0���.'2C��u�iUm"G���'{+�G,�K|o��'�њƇ;O�B�*���^��.�K�16&�"J�����z`4��I:j�����B����+��ϥ���T��\䧲R���J>�]Kg���jL��c�a T�k���jq���m�!�!k
��`VB�t������}��WSm˧F}wn�W�JE>��D-��琇��C��Q�M��*�{���gN�o����q$��X�Ͷ�}D<	�L�g_up*m�tsٙIk��Ɲ�R ��D�Oj��}y��g���ڍ��rM�}���Ff~*�^M}��f ��͜'��fl��f��/��$ƭ�r3���z�9L�W�7U�IN�S^��6�A�XRv���n�4��[T�VCs�M��P�:�$rM�;�Qa:Y�i���%���s�����Z�hѧMwW�^�{7ؒ��j�����-�R�����?W�+s������5;q����[�{aV���PZpҼs%��[L܅**�Y���9q�y<���/�d"-	�����O.���	����xm�Ot�w�)#�и
�F����W�SK~v<Ý���I����s����~'�4� ׼��ϋ���;����-}�x�"�$u>I<��d,{��C��-��%�ܤ�\l��%?MD�׊Q��B��Q�t����Χ_�#�=Mk�vrC���g��\O�3��#K�������;����U/R�m���=�a�L<���1|_�H����{���)�c���fr5�e������'�=%N�~�_? U^��S�8\� �km&m��,V��x��)Ԕ^H�x)W�����;n����v];�<���L'�M����'h��~%�!��͹�~��Ԫ��y'Z���y�*��M�M�������h���VT�RQ�f$�T�~ˬ��w�����VQ����x��5`3������|H���V5�yhѮ_�>�|O[r���5%M��g����r�M)����IE<$���8-��Q�˘p'��}��-�7�SM,�(���,J��A����4���|	�i6)��5 ��\��+.v7���x`����@����SZ�w�i��.;��%������u�n���[���?��R��#��Ĭ�8cӰ�t����2-�"�.aQ�V��Җ�Ѷ��׽3�T��y/��c�V�y��{�L��f������ZX�/���`�4�и�x0�fKJ(�<'�Pc�A�3���6���/T{���u�����_��*1�r�f�/�?4������S��^��Y|���ֽ�Z3�駍R��������S���~�����t贁����?�'��x�����IQn��$�s˸g똜�`j_�iP�j�������?7Tu��\�y9����4Ī{�x�3�߾F�����[DYf5��ҺŁ~�\����P����t[�����7yTSiq$���(����?zR��Ս-��:��ђ���+��E}�˰�	[+�6k���n�fKg!�y|�U0�z}�����g����=�N��UmsL�w8����<|����܈��Cǖ+�i��W,|Sy?R��!�7�bZMv�|�׏Q^?���b^�D(<�6�a��nFKx��/�H�͵iryX�:*��G wu₍q�a�~����\��3	`���hr��Z������ƺ��[{c�z���V�0�W.���p��fRi�4~�#R?��zhĳ3��n#�6����[���Q��U��n�$���JK��@BY���0i�2ZX�.Iq�L��� Fw'ݯA�I��xZa����S��yvEE��=���K�	����%/-�Ss���R�;BTC	d��l�+�U�7���C�cuӜ_�Ϙ��c}���r��+���k���a=PxT�|��a	O���Փr�:��cs0u�&�Bס��~䄟������k���T�̫�n�̇r��ڒX,w~���yj������H�
�No���M2�����{s聅�#`�Jsx$ߚ��{��Я��/[����]��;s*��p�[�v@���ǎ05%֦�q�i%]<~x���߳E)�2�L�O�TMW���D�J��^0��J�����l�+�M�]:�,(*Z�§� CM��qo,���E_%8��N��֦w�U�M�g��s��4u��K+�����wo������f�$4A�94l�����N}�
��fn6ƅ�\�2:QV0�}���Xb�6�}�ɪ�9S�3�?b���^��JS���k���ORs�?Z~�[�s��1�C��*+I_7�	wn�Z7�	�bMZM��y�z�����!�z�,�v��|1��45�Ā��P�ˆ��9�n�Kq���񝥼ü���55/3s��f	�~����X$��?�Z��c0tZ$܇�(�'�UUF�%�I���v�\��9�H������I���Ҩ?�W=�8���r3���2� vq�!.^|yCFޭ]x=n9h>8�5���#dk�\�&wfKڮH�j
�ZzW�#�.&�=$Q��m�����cѪ5�^�:S�Ʒ���ݛ�]��[_1^�n,z���_�L�w�	�D�����~�LMI�Y��2�N�sn1�92WY���h�̔�
���S�
����p���UUcqQ�҂���&���ɪ���9l�����P�s� ��_�j>�����8D͉X-���c�f>��Z-�Ч����G�١�)����Zy��E�f��!��>A\q��4Yp!����r{z°�-��[�P�q=�N�d��i�$��^��p�B��Q��D'XY��8G&|9���{��n��f�M�P��;���k,�\��j(G����<n��G�;m���ld��`�lzo,�Z������$��a���j�qu�������l��}ޑށ��Cφ�~~��x�:U�^�=���C> fO�p��@?\H�/��K�;���T���5��,��V�V_���s��ijv	��ı�y�˷2�V�9���ē�4YR��r�& qd�U-�X񼑠��b�Fi胧�|%��@�������s-���y`�v��}��,��.��݁*`�$�Ph��~2�դ`H�'I���!Y�Z�/B��?���$�P����>��\ʽ̸O@��O���[UX�q��@x�1r�Ou�Wc���4:z��l�ăK�[�9Fq�&([���������֫*��|�7��~� �U�8�դE��\���i%_2^3�(�m��߷�8K�XI�O�����ݤ�z�N(`_�e}c"b�o��7�o���,�
?߫��1�+�^`��b�	9�M��F7��M�'v�^6A�=ʿ.�b%����>j�5�>�蚆gx:$5t�$���U���(@��?�n�~�t�\;Q4HK�lev��E��i��f��87�->)Gz�J�M\��������mO�@��mSk��`4���յ��l��/D��8��p`����z. �7�ʫ(p���}��݈���W���޻����&-�r .�q?$�;Z�>	�~9�jF�.s��[ӕё�޿:���//r�=	��pO��`8{�r|�ZnΧ�xc����'��ػ��1ڪ���n\	��
W����	��Gtp��`�o�",,[�����Bm�5W#�N��HNӓ�F���K@��F<�N��x뮒lK��]��0��OQ�����a4e�2�� Yc�/�;�{�?J����pY���3)C�����9��S�Knf���<@U���Z]t������;J2^'qR���*b	U�|���A���d����ӭ�쳵D!�!{iN��G��Ib�.V�r{� ɳ�S(j�=p���s��י����+�}�(�C�ʨ��Q��9�Mϋ�s�����&�]��f�F����n�8y�s���;���9���[�y#_����˦w�83���Y�Hj�����HU9���Q�)�����(��X�u?���5��1N�>�y������I����9�T��9�j�[q�n�iI�'X���aS��I�@ف�*ǕW�2Z���JΠ���ݲn�t7����M�O�%�w���U���5f^;V��3>2��!���A�9,�u�v�\�q��F��Q�V�ҷ����6�Q�5|F�Pv@��3�i�Ⲏ%z�2Y]2��F�͒?%hB[�1��	�̟�/(���oɺ��+<w(.)�|��|��V�����G\+&d�p
qh+����������a�s�b��.8�m7����aX�<�r}9$�j��ŴE��b��G�|�b���e�=�H�C�3������%|z7�so����� �d�Sޗck�g��S���%�Jn̴`6{㘏dD��+��^m�g�����Q\��x�Dў�oK5����]-���jX��	->�y�Z��2��ƹ��\!��P �'�*��]�����*��f�_��)}�~���ߙO��&U'd5ELązO$f\�	��ʭt�³��]����o��#�z�n6N'������o�H(P����.�wUqm�4Y
����#�־O�p)�������L�sGl� �&���$w~�;�Ζ��gE3��I����.�=����q�0���4��%��UE��6�j��Rh%�q���2�c���D��P�(��Q�n�K�g�D��S�B�z&���Q��/5Q���ۋ[J�v=;9Wa�9�����Xn�*&+�֯�O�٫��b�ۤ�ȕJ�Q��X���;�LxQd�7Ђhs5��my��r4�C��̳�pwDS���ì�)����I�s��u�d.�ܰ�͟�{!W�A�U���^����e1�	/���#F�֨�)Q�i��G�6�8�1�9Vcj�]u���>{QTl{^'������J�9/��d�I� %#�Vw�܍���JU�V�B�ew�Z��c��<�+f��p%dLz���j��ar{�-�]��ofK-o��Sl�lܢt�d�45���/�O�W�O~�G~�}}��	���jx�R�q�]���|�
���ei!����N�߭M����d��@c����v���>r���b��~\��-��A]_���F� ���o�euA�i�J���
T0>ُ�D�~�ևO��_/g,�~!�V�0=iL"�iG�>��F�	�L��g�#4k�biDb�xn�g�!.ӡ]&�5Qa����2��K+�WSm?Gl�����&@�3a�� 嘶:ljwTZfqf�bJ��ܱՒڿ��5G�\�ٱbp�H��G���ˎ����K����MJMU��b�0+n�Ԡ��wM�4t�5����Ծ��X�7a��aLt;������>9���V�#,�!�A��8a�rqJT^�|49.ͅkeaw�X0.$-��-W�m]�X||�ւ!I���?p)��j�_}��}��M�Ms����K1o����n,�Ed�j�}`T[�Yg��\��Q|����NL�N�o����[6�gʫq���Gu"��U��(.��ʜ!L�zC��u��vx�uڲ��X��u¦�����6rӬ��� ��}�?���D�V!!)\�/�I���Q�zZ�K��I
��_�9���&ǟL@�x~�O�����T"�W�]I�c�zW�Z��P��������їT����-h]+���T/L?|+LM��AW�GسW�o�����Hc�Y�ʞ����a�|�</��ۧ�50²�(o�����u�dk,�#[C!������ `�S�Q�g1�U�&�6­;��O�k�C_&����Do���"���-��a�ːx.��v���o���hhwq�d妾�g��T���7.��Aܥ�<���k��k�㩨��puRӘ4��Y�#ɸz��ʃ.�Rr�R���������d���$��'U>;j[|9��J����dP5����i/|�OF���)�=� ���K��X��[���2H�;}0���W �>��4�G�Y��Wf.Qذ���M�r��٭�8^1(����;�Q>�֑~z�] ��v�qW�}�`�Z_-���Z7c�����P?��mFP�Y���xΒ����]s8b���3S�E�s�x�F�Bt[Hu�nF�W���q���"�1�ހ.��	�׮I�6�wn{��8�ޱ9�(�;�
�g���B|n�H��x�3T�,RWk�v�	�i�����?;��N:����*���	B-^�&j����<3@œ����'�<ͧ��}j��!M�7�r�:��D��j�2�n�?[ĝ'_��8��h9Wdr6�lj�-ݺg�L����F��)턲R����
7����?�m݇Bk��05�1rԡ}�	C�
���t��È�k��L��(���Ro4��&!&�8V+�:N��a��#$]��9�v��>��/�����(���c��u�?�Ӷ�ڤ�|�jb�>tE��'G���}1ۚ�i=A���2����MM�{Q"���M��b�˥�kDO�tʣQ�Ζޡ���Q��䍍r²�z�ګSӸ]�j�����CA0��
����x���S�?j�=k7��<��V�	��Liu�*�V��*
�]�g��O$)%%��.�s(��ݓAH��]0�$�>PR�$�������=:��������"�޶�[s8�G���Z�RU�IS�8��7�F��8�2�̬U�;K�9x�L����`�18�Ly���~ΐfr܊�[oݿ\����I���1Ae�����?�<���}�ё[�q���>��E���wkZ�9{�������S��P�L�B�y���Qֲ�=�FG�犅c9Q.�i���d����κ�MI����%j}8)��q�C��6֕?g)�G6�O�zg�ȗ�XN�MC<����b��L�d5���Ё�+��_�#�YokV�w��[\2���U(�fKcJ���G�n�Oo�P�6��
�QS�\0��Q��Ŗ8Z'f)�̡���>w��@'����S:�՝���C�l_�C�u[�8�sj,<뼲t��@���"�jio	��$Lv����uX_�X܉��<w`�X�򿏃�o�(jhP��M_u�����?�s4�f�`����\�$�P���W�[��֮�T���((�`+�e��r�3H��,�6�6iZ���ěU#cb�s��,[`Q���k�Hk^�8���ͥ"Jٟ,D�r�՚'@�Pl��8io.z�ѵ!%���$4��/�/��]���������,��`�s�.��L�[[��	�o���=0���dƻ��S�1�1�r(*z�J����qJ�B��ʷUD	��Yӟ��G�d�� רy{pv�r%I_߰�DaQQ�4����
Ԑ171˦�y����>'��CQ�T?����P?��[-���ݞ�J׉�n3�N?ޚ���X���ܸ$_�Q��61v���k,�ݚ�ӂ��x����k�#��o`S����g� xG�����b5���O5�Ʒ4��9N�rRb���nJ�\M�O���늑��5ϲ�ػ����� $M~b�*QN-�����\x��64,��Z����ݥ	�#�y�]��v�>�k� ���ΰ��3�v4/�L�g�=CƵ�h���D�H����N�x+F�-�2&��%O�c�ʅ���s��c��ZQ�{_
����z�e��}�ݗ8r�=9�:��4���ϧ�ͳ���m��t���5?��)�Hk���|N�>r|���!��,�]A���<Ә���ᚤB;OP��>����m���'�.���m�8�EY�$ޫ�^f�y�#[��u��\��S������&Q����f}��U�\��&��ʭI3]�f��(�j@�L�I�U��WP���)�C��P%J���QI��\] �ã�"��N	��m�G�dX���׎6tJ���PpUC3�?E��Wf�����7?��i?U�i�|�z^~���(���n<_���>J��5�w�.i� ���d����G1G3�!FK�H�a�6�>7���pA�DvY'wb�G���_�Wc���##,
�?�D��7 �H�'��i�p7@y�K���"{�`R�ؕ[@o�Ժ�̦��+�8�!��R&ܞ��~k,XZ=ן�F�+������z9���n��T��/ۙ��ԙ�!a�ݵ��)|��a��hAv�����Y��N�;|�;�A�!����0%��sё�Gh�/�����R�7�Ҍ��ԉy~��v6u*���X�^��8������M�y��`d�p�;��&Y2�&�S�z���%�[�~w��x����ܩSuL��7��*�����!�@�wX���Ӳ�!#�~�Dʻ��ɀCTxJ�VS�3���pa��c9�2����n�l� TUQ�RE�o�.��(Y���G.}�?�<?�ɜw�����%��q0�8��ѯ��G�ڷ؃�$�r�=ޚ)X1��?��ϭ`�gX�}�V��D�����yf��-3�\�e),��c�|��~��;���J3�yMS���4�@��&�*���"}��辟�+���2	3D���p:{!o}�-TT�p��$�45���iş|�qذ�3�.s���V���[2��tzj�T���S�v�)2���A�mPc���@�չ�\Uޮ3�ey ��� eŕ�L�yJ;���Ӽʃ=w��7�s�+�¯�R�T#��&����b�n��4��,x�H�w<�n0a҈q��ֹ��(+��w���u'�T��o?�V�9K*� �r I"��(�F��4?��m����9��׮A �U]=g���$�3��H2���뤢4���#�[����`X��}t���B���\�H�#��m'>��ǭ� �B��/������#��Z��MU�e�D��_��^�,妋�X��n�H3G��<��H+�]�oU��DQ,24K��� 3�}E
��R�������L��uxز��,�:�c_��&��u�`f�;�w>�TH��4�	������:�d�~f�,<U�Y.���A�l�k�[��m�����+�9�#z^F`�OJ�:E�nf+}�G�����Pe=;��|��6�Ճ�.jf�A�XSf��'ce�Y�Nе�.�龱��$��\:)&i��Ӽ ��#�ӧ������Yr;l@�kzz�+�σ\�W�x�j�� �V�S�vs�8�z��y�d�#;����54����Q#�.�Q�)����߷L�L��m��!�(��\'S�Z;��5Q�y�4 �3e�H��u9����"�2v.���4⃟��zaʔ.�O\!��0�֫]�rL�6(�~i�Q���\�P���20̰����J�|��즺jc֕۞�{�AR��G�ϖ��9���s�wU���ۃ���-"�턀���"��m����'�JӋ�C�s*��{�^�<�f �����6:|��Fl���k���Q�!��K�]q�7�ub�a֬��4��|0b3>�fb]xd�l���fP���d}�H��T��`�!1��h�0%~lp�)�F��m���G�̮qE�����\�h�tbK&��ZP-������zǞp�r�?����5~��I�$���r[�[ǘ���Y���GV&儢:d��XV*��Ǵ�����D����Kf���4Z�z�	*$�?�<Q��uh��d���rЪ��KYy�D��7K���6����ؼ^�{C��}�c0�xY�io=,:X��X�һv��iK�7F4l�]���z�lrf��TG	�뮭������g����8����Ô�ӧ\p����$hms$�I����R�t�]�СI�d�ҽ�� HH������e��b�KQ�Ј[W;��U�ܥ�S��b?���t�j֔�&o��#{�j"�%"h��A�_lR�ΑF�{&{چ<�����1�z��Yw��X�Wex)�X������ov���|�UK#��!�4�:��Q}��L�% Ŝ�.���s�Ŗ|�-)z&�7a&+����X|����怬�G�%β�/��.ƍ$���NI:t�*־:Ww6K��}��\t�X����?�����3�ڿ�����{U�����e���!�,;��T �x���e�]ͬں����s���B�wΌ�צ{��c�t�/'3!�<�E��� и��z�����$c�C�(�D�1�K��~���T�q�jb�0���D�[s��V˙އ���[��8�`���B����j����Vu��:O����t��c5G47�H�f�pp���;�&�>����V��i�բ�@ا��ޕt��" ���K4���V�Gޓמ�?��z�`��k��~��7���]���^�
<���|�_L%)��/���Ε�	w��ps���Pߖ͐�W]���{���<Z�k�16�����\I�A��Ղ�b���G6BN,������K�{#;;���ǰel����j�fA�xi���\�qN5D��������H���L��_N?x8��}�3~����0�>�&���	�}��� ~[o/�����Wm��������
S��T<A��̫ip�U���J2^�V{AfKm�} ԗ�B��'���7�B]R�������L�w-<o�1������I{��+ħ,1�&j�.���pA��a����Z2އ�,�_-'�5W�F5;���U�)g�eNI�Z��՟��|�k
�*P��c��hxO��Bpm"g�����>�jSPS`�W�O2h���|%&��\�Bw��]26�_{w�!�q�B� �0���!E_oΕ}.�9�˝���Ț|ay?Tr�6Ny�_i�R��=[�t�(�Ec�il¶�>��u��� C����B��� ��ϝu|�/�}�c ��X��y�
��U�������+���$'�H�g�7�g��C�&�a׮��*�2�py~ �QM���q��GC��nU�F.�Gg������Kt��/k|mA��4��FDTG�oX����4�3��M��+n2����k�̏?�Ȟ*`������^d}�i���1�v��+��G��8���m�6�CL�)���y|��Ȳ��5���2&^j7ם��)07a"�+˒<l�����`���w�PK'ٱLÖ+eO��)[���US�+�c���b+zA�&��m-]��9��"~�ӗ������vv��"��
�� ��2�1��J?JC��'��(�-�oDC:E�D*$���ʠ�*�r3@��?��Q�>��;�A$]�>�v�mRy��/�`h6z	�_�|Zv}x}�,z6���Y�)�E�lJ��'M���x#��e��,r�|���eg8�v���n�X�����K��5C���{��E�v2�G^#&�_�<�)-�oX���1�+1H��po��(���ti��+Rߡ�D�u$J~��z�P�7��O�Vp��%�M��c\t��>�m���Ԝ6d�Z��ˌy�����_�7γ�c�'D�_QJ�,� M0K5$0��,�L�U��.�z�$�N��3�Ù_�G����^|p�џ�|��;T�C��Y9D�<$qa���h-���{��\-e��)�i��_ݣ�"��N�^^>	��."��4��^�$�-��٣�EE/Y��~V�X�G��1�H=�L���m��9nؼ��F�d�t���X���c!�#A�W�~��xy�������HŶ�u���<�D/7�Z�ф��T4��ę&i϶�~T�
;�4:?���:e��+`�<�WC�!L]o����!!6�m����`Ǆ~
��|��X��]��y�7LBm0E���)@#H��v����Ԙ��S�=k�Ұ�Y�J��j*�E�[�Ó)�+��MkZV^a�-�=��n�����_D�t-���ߑ�ٍ�$;
�`�7���d�/�?��||�4Y?��&$c[I���vwcJ�*挿�}U?c�gF0�<��J)dNC�Zr��_��$�o��R�<���y����[���I69C'_r�M�np8����MDUk�[��d�E���GOܭ��?�6�-��t[��[_?:��� q���,��c�]/���Y�_�:�ƫ������[���6J\�k:x��ᣔ�R�~������"�廚���ڽM��F��A��q�*�����R����6L�B�A���Ɏ����Y��@�3�{�e�:�Ĥ������w��ϵ�&b���CvS�J	�h�f�(F����syy����4y��2�i��'5�
�Eϛ����:������h���ʨ�Q��ԤC$VS�瘾����
[F8C	��"ϻG:��[҈�������^Ɖ�N�V_I8��5_�(:��n������Ě�l�DW[�.�~��m�z����S;4O��t(�(��)��E��e�7���ؽ�ٝWjߢ�$&���:�\�?TTU����ɳ,取p���<;T߽d������3W9i!���8�t>�h���h�Z�����|�� bK�x3�u.��qл��[-x�]JT����AA^�G������A�����!͔
"ª���rO���g�;]���Tۖ��|�x^�k��o��v� �?~��[ڡQ�q+�.T8��8\;��_�P���A<C�a@N�x��0�ĚhUwz(bW?�҉"���i`�񃚎4�`����o'�K,�٘�L��ᒸ��+��@�y���]��7Gz�1��'[S�L`�{���:�G��P�u�҄vt.g-����ʘ��	�����zPdC ��~�0�-�k;z�,�IH�xoٳ��E�Ƞ��ez����b�������G�K���H�*c�ɒ�tk݈A��:�����G�Y�
i�95*Vp�n"@�K-���!�۶�Eڏ\m��ݚ>�v8ZA���<��<�Ѧ�]a��Wӑ\�.��I�m�����n��'W��xH�
�v�<Ү�@PM�S����T��`ʻu$�}�C?^�Ry�b�`�]�;���@�FS��dSn����#�{�).͕���.�p8t�~�[�K�@�������7����ʻv���^�yA j`��W��65��;S��$�1�Kp���2��"����n����a�v�^U��ȱLث<-���y�c���e�V�xΨ;>�h�����șp�uA�w"�&�dJڂ0�S�xi����j��O8.r������]�`��ҁ��G�������v*������>�s�m��,��n���`��8�Ӫ�;!,(�Sd��@�
�F����<W�s&R�1d�`+��n��� ;�����q�QQ_�(�%݈JHw%� )�]1Hw�����-5t	��9t*͐��s��������ݼ��=��O���Ve8�HH)�7s/s��ܨq���{,�]�*�����&'kh�V���3�&RY�6�]|ݣ)�Vh�GXٕ!���6����)I��c-3	��a�,�e!n�!��M�y%8��&����'���)	����7���a��b�������\�/k] �WA�n���O����ក^K��߲�����'�)=��)RfD$���޴��̛�9��u�]cX9sS8�},��;�R��7��Ơuh��Z{0�H���!2{c���z5�����t ei�M�K����mC���0I�=tq���.T�p�H��L�a�B��ke�[���W=4��2�:���70H�pg��bP��ecL�)�l�e&��ܭ�8��8�Ȳ:Z����WT��K�=;�� G������i$�3��W�wu�9=�I��3���=�*U������ ���>TU��3��li��#�+1����?����u�"ת���r��(e�*�{6Ș���d�[��W�WH$��=:i�U0w�İrh���8�ޱ-x�oK��+$'�����E8�֌����P]iXظ>�WjF�>&ænq�ye���U��W�g�|�*ݣ-���� �^�����_yu��6X��Ѻ-������	X��Ǐ������+2x�F�������aYz�滍N\:��/ �眈��J�m�c@^���>� �z�E\�����R�K�A)*2��"j��y]�W�(�����/��K�+�X��3��J�����~�EҚ�7ؽ���g�\���=V�!\�	|�NP��I��CN��_�Í6k�G�ƾdc~4n�ֵ����b�����Ї��`�o�(5�q��ׯ��*�+F_����=V���=>Q�e�Ɋ��Q�Q��6]��Β���y��w���_y��N�(�U�ɔ��m�;p\��1�!��a�b��4��1	g�^Ƅ���������9ù�(��S�Jx&c��"d�G��8_���o�B.�c0Z��,K������t�D]*�K�?���{���P�M;�eİY���5SaM���%M����F��?��~���ށ�8�on(a�M��\��v1�N�CGUe��}�H��Qs�� �NP7�RId h�l~N3vO��Y����q	���M��#x;u�0�
R��:��2ӟS���:ϓʹ��������e$l��t���;b���z�x��;!��pA�7��d����WcE7޿���������"�XO�8��D4c����RW�٤�y�E7��J��!F�u�=�!öQ�n��⚂�. �h�C��H9���G��=?ʇU�.Zl����E�U�N=�Ŕ�z'wy� ���jGR�F!�h�D�etF{�י��Đa�(Ϣ�@��}z��@�:LǦh~X�\�xy;�be�o��觏���80�0�V��J���ڣ�������;�+����h�t��G�h��P8g�|Hhu8�����)?�L�\��9١�;�(���IM�oK��͵�n�lɲ,n�;h�w��� tޒ],����LHh�>m#��u�.ueJ�;���l�A�������@A��C�z��IZ���V�9��
�GkF1)�,,�"3>>�1@�?2�4�f�k1k�2_���u7עҫ����,nX�����[fpsN���S���3u��8\"s����_I�����c��O������5��c.: (���V�&z���C�Q���R�WIj�(�k�����I.�ޮى	u�8��d�><a����<T��g�Ϯ\��;��%�k�ʶ��=D�i��2J�����eK1udB1�`)�n��4U�2�ۗ�G�$3�Y]A��Ÿ�^l=y�i��E��UtȲ�� Th���V*����8��Q����1F���kC\�G�5o$�oQ�W�m���S<��~B�85�|e�B>��?D��N̬u $|�v�G萇�^��l��gc��J���d��ҡ��W������ٕ�E���n���[����ã�R��b��o"oB������WZZ��Ŧz����}�]=���[���j�Ƥ��� ��<����]%-~�ܥ#�G�u.*��q�uT�:#�_���cc1�Y|���4e�g������Sa���43�R�/��Rn�c0�K����˝�lwPkc"J\{p��uFx��Y��]���e+Z͸-�ؔ 	�4�	ƭD�b������[	a+�wd�n�]�$hX��e��f�SS�_u}?J'�@���u��v�h��T���<a0mеĵ]f�H��V���'����\ߙ��4U�_i�sCG{�B��w��N/kT؞u#\Qd�?9��UJE�W�_&x��:����zYm���P�'��n��	u������09��E�5��铎��[}�������V��Y�����8�]�_�0wv�R�v��@��EE{��z��k��x+�sg|jZ�*6����ᘇ/l�11���G���
yfr����R+�j_�.�|I��g]�3�2<8����g��[,��d��*�uV3!����h���A
L��*�X��u���څ�Ra��=�n|rGQ��(߱ٔ�j��0RC)q�����r(ݏX韫��wT���.�1>GG�9�AxIW/�[�D���� /�z%&BJ�����;�`��_��
0��l�]�s�N�(Y,U��4�,�ι�t��[{a�д��[�����!���)�C����\S�~��@:�i� q��vk��}����di��y�5)��X��k��:Wmċ�Ӟ����������-[Phi��+�eb�7h|����t�L]����N��T�$�۪�-����Б!�2��Di�O��I�Sl�ޢ�W�������ՊӬC�ɂ�L�Y
k"�/�DA���_�L�p��#���&��|�Z&/���q�1D
t/�d4�A<]ƣ_��+ܧ��J��m,���ђ�-}(B��"��\#�z�~���3�������ڮ��륍ol7���'u����1���ֺ�J�Su���, ���>�� ���dĘ�7=��a�޸���5ʮl���*�G���.�6�ő�fҰ�{�����>���qK�� o��@zko�~�v(wCh�v�f�u
l ��Z�k9s�6���3*}�s!�X�� ����Tݕ%t�LTUO�lpc�#���mZ^�,[�k�����vQ/E�8�o�� h1�1�O�g��[�}]Y|'�&��_���D���u�PT��y�0�)�c�2Ԋj��m�^��!sGi�Ǚ�^�Q�k��Q�Q�����(��rI�o���>'�?n��=���-z���gn�% �&����K�	���	�7(|�`<�GcRȝ����#(~�hFS�ʇbj�x�Bd�k=p=�ʩ�=k�i�ca��Gi���_�����jM�[m��b�)y��F:͎�����﯉KwM\y�i�L��h�;<cs���F����t���,daV!�<k�jC�_��n!��0Ӗ/I���ݘC��W�\
M���]e)��cY��-0,O�xw��X"�m��Ξtk��9�}8�k�u�B2>��y�s2e��e����К�p�?�(�.) �[�"��V(�r�C�;с���+Gw�b�f��o�@I�����P�H!�B��Lst�o:�,O�=�mk���jx#����U�����]=�V�u�g�WF��[vN�{^ɊL'�W��.�H/�]|r&���3����AK[�o!Ww}m|گ5�t�T�`��PT�0gU�H'�S��~VM���J6� 3gl�սP��ז�_[��گ�:%��mG�pP�5,0	Iȧ���f���$���>1�m-�a��)	��4�;���'	��.f�Ɔܞ����Z�#���V��i\�;zyy��o)ڳC�T��p�6�>ǐ��d���L�Ѣ�J��*�$�Mٛ�MY)�]����r{a�B��}���P�V≔�1c�c�{��;���n�ˣ���s�^���j�<�T�������Q}��4 ��*�m_�ǹ�5_�����M� �4٭�'/Kt�.�3�X	�r�U�{�z�w�R�z_S4]E�=hn�����f�i��h��ʈ������������}�ٸ)�C��F9ҴD;�F}|s�c3���g�������ق:gz�v����fQ�7 +s��~���{(���xX�+d4�v����cH�&6����1�1O�f$�$Ԛ:�����˜�D�u��o���z���m��5o}�f�C:�^�a�� �=���XTN�~	�Whe>XS8� �7��,N�юۚ;��|֏IJ�2N�b��,8�~Mֳ�+��Z��b3��Y�Qg�E�w���G���?��<���.�n�6[�R*��`٫�dV�8�H�//�T!�"t5�>^��8�Ԁ���m���
�����7�+���w����͚���S�p�E��Ҵ�@#XYI�b0�ã͢���}����jw
ٙ��?���2�3z!(-�q�t�Z)��M	DB(#���܁�ԃu�c��[�{��tB]��wAނ3s^2j4#^S�qB~W?`���9�5��� �3G��������;,�-UK�9�����Z�ͅ�%!� ��E����~���Ͳ.V-;��ҩ�X���۞U�K�KҘ�_:xZ;u֎Na�c��0��'A��VW�@�0AF1��q�{�h��
�������׶�[��s�g>F�?r�8l>p�Fr�	�r!�n��/k�bw|_k����*�QV�P�
]��0��$�K�t�� ��w��-�Ks���ɪa~�g�u�P���:Af�7��f��'����������uQNV��_
G7��$4��%n���y&,�ܚ'�ICNrP���+<��'���=tH	z��j9)�{�O����e)�u�j��Nz+mxLҹ���@���ر�C�W���I��%��|��g���l�Wz������+zN�[�a%�J~��č�a�D�,��<B���������)^\���RC>�K���%c��S�z�Q��c@H����� t��� ���M���# ���������DW��Ѵַ���:wt��E��m����3Z�.����G6�^��~�<��e����r�6�<o+'%G�<5t.E5Y�������g���Ȅ׾x�j�@����]�����Ł>�=i�ũ�ܼ~�=V�(R����UM�B��2������&��N�ß�Ph�����V�&�>�>��W��gt'҅��C|���
���1���&/�P��Z���НI����l2B�N��{��b����@�Yr9~�]>�)������?�^��l�/.]�*���e;�e8���ke��|Y��nf�3���i�T�K�m5����&���Uʶ��W�1:��E��-u�FM������]��~�
��fO{_��S��t;ܞic-��T�G�$F�%�i�54�JWY9:��~u>�+�	����h���aBE8����0	�ġ��.��4*{��I�3)�:���\mc�8�$�T\��S��SY�Ni����Y������=�|�ڞ�	�D)+���ߙ/�9v�O�Df���j�Wv�4§̷c�d�,^S1ݤ�~�`m�W��iWg:k���S����b�.��$E_��;U���Mc@O9��
�*3�\�s�gL����R�mPI��
.�'�VP㹘������j�m����;t��������ʶ*�7��3S�쿝̽��4<��������00�z�uw��Ĭ|�/�,�o�(���:+)�&�νH�u��Xb�W�ok���r@�t�����!-�`/�o��()�wq;̕D���z:����?�h9�+T����j�3�!���RY*�_��m��J�2]2!���}�L�X��Jߟ�9�g	�Jvեb#Z�-6��P�DL; j���[W��Υ�����G��ȵ��Z7�{�O+��e�M�������YVאw�L <z�/^�� �pe@bs�x3�_���xR���}��ܛ�;�Ҷ��vh�$�xg䇭�@0�^��y���>셈�y?�k������s��z=�r�����*.��5�kuZ�gY>0����b,3�h2��,nywW��x�e
TrK���S��8ͱ�:jO��3����ԩ�H��Yq�$�E�vCF^ұ%0�eS ߦ@%����5.2���2ED�{?��#Kh�5���t�oj2-OU"���{aQ�,�cB�+ӹ�7�'�C�Ye��[������}�����&���-g��݋u�'���_�.�z"��T�+�n[�ҧ�Tɣ�#�Um{`���[�� Yه}�P_�e�K�M�e��q���4WZ�ii��b�ɖ��C~���]�9r<��:e�+��
3����R�F� R4�ߙx"jHf��ETi�.kD��E�:��`-7��.���}�rbl�F�yN=��{)ۻ(TL6U�l���j�[�ļ~�)ߕ�8��F�gw�1�=	ΜB �պ���q�G�%��C8{��q�^�G��V�A�%�ϭb����S�f�^�E9)�UKևɇ���Q�����8V���-3ƫ�A�����r��y{��-��S��W�p�MT}lW;�	��һ�"��xOI$:���tq��!����w��X�i4��-o�zef`�:Y�mT�V�kev�jk�\d��O�d�eј�	��Z�5ze���^,�^A\ev,͸w=yL���X��CƠ߇,k�H�(e
K������=̲�d� I�<��#ϸ��?�	,Ӏ�͌n�\c[����H�Ds�ڨf��^�b����F���Z�����r�� ���zK�W���,��	��8�hTT}�Y���I�z;���
	��k�&u����Ĩ��Ʊ{շ��]���*|˥���!֘q��&�����MӋ�.���~2������ĩ��

��̥H�*i�ш����ܐ�e�go���>De�T��|j>:n��$�����E��M
�����9���(��P�w�$�#��jF9r`[|�f)�"���H������nGd���AZd���X���m؇�Y~.m17ܬ�k>�.�PB�sU}.:(�[��s�3@��.;�i��b�W�#�$rh������P-�BW.N�'�4_��C ��Z��U{�Y�ؤ�M(�\ �l&��%��V��Y��	4�сޱY΋���ʧ��3�ɐ����%a�w�ɓXr��q�Ԙ2;�t#���;�d�{�f<L)��@���"`ve���5xk	&E[>Qh)+vHs飭�gYږ#�qg��i�WH�&KC�<�����Z�vN����ߜȌj��9��M�4p;&�W9g��n�����\5�۱f%���`�!i��G����
�L�����I��̤\��lM��Y��H9��z[!߰�o���K0H2P+M{��A���Q��\ߘ��($���r�!�+0Z�;ʭpw�S!�Oq:��2pSe��#��j_��.�odF��x���X�ZD���t���W�(HeD�|ޛ��̉1���&�l��L��ʸ���	\;�X�d��ĵ�_=ު�c7)1�.�?t0��.V�P�X�O��n/,(�����n]p�K�Z1a���V���ǭ�����Yp���T����b����}[��C��!�p����m�ml�za���׸���Ix�|�+8HvZ�{�q͘�
C�w�h.�t�[���f\�9`���.˶���r�D'��9�5�Yn�8�{���;"w^���-�O��='�?a��;\ڥ�Jo����#Z�>���p5�����jG��53��P�գ�"�6�po�N�h���6_��]Ƃ]����!2֜N}m�ﱜJ����zy4��g�\�;�����Le���/�����M<K��L�:4���>��o,?3۪�/��5��4߇�U a��'X5e�g޹�"���IET�ÛdQ'����J_����ir� ?�fX�wE)��cc�7H�f�CI�7sXZ��c���)����Ne������$��#�l.��f�趫�!��?���7�H�� ��F����>.�^���TI�"����3nh�M� +5Qu=��o�7v��b��n�\�N�8��>��^�$������:8<���yZ0�U`��P���[�`~/²�{��&춅�q��][�\ ���42�u2�=����)�>������J팗ĵ�٫�¿�B!w KL/��*������i/�{��l��K�~Ԅݹt���K�v�6ag��}B��Uݣ1!u`���/G>������!��⠡��2� �&�	8�;8�gf-?��!2�G��A���)��yk�-1�5��pR+Wg=ic��;D/�ܑ������1>ӍG�
$0��oU���5�E��6�Ƃҽ�k���x�g�����I@�3t$�K^�����F`��/]�6YҕQ��,��*�+Q��Z�\;/?���ޓ�%��V��$�7E��f�U�w�~�eM�(!���f)����h��v3k��;�"���VI9:ֈz'��'�ft�L=X�� �G��G1j�KH��k�'�"�\L�QEyw��YӍ�h��'h���e��o����?��N�4~�|�F}2��v�kGl��hs�	���d:�&ŮfA!|�%F�S�� 	m�x����z��ɑʠ9���_ȼ�[�:���/��{CL��z-�M`��QE����k{�E��o��X�:L�O�9vYz�7?��h�yř*e�W��G&�7b�QN;;�ؘ��)��}�������� V�-�����F�G��R���n���Mf�0D��6�K�����(�}��'gm�&�[�6Uѳ���&����q=��{!�QR{>d���y��PT�}#�T�����oZvJ>�+����݃�9���Od���'�f�w1��L|/�Ȝ�:�ùFO���J։yYa^��o�3�_i[[�E��ڽE�/�J��G�Ji�+xmKu��GC�z�9�H�Zy>��"N�N�mQ�fmm�6N�V�i�I�u�zi�Ǉ��3��(��/&v0^��gŎU8=�����>�B�م�	'�x>�_���?���}-;���N����hQ��yެW�3�ֹF zX��h��M�?�ħ�%l��ڡ��-#b��^%��U��Ws|�=�)�^���S�����8�85�\��O�Usj*#9o}��H����kX7Eo�}GW�x�l�˝)������h��������l��}xg��z���9���QyAĥ��	~�7���߭�O��N�W���5q%��|��u�n"�/K�
�ok�:��|�u�m���2���� D��Ϥ��6M��jh��/�<P%����^9�+��t�����e��۝oz� o�R�TI;����a-9j�6SƽX� YpЮ`���5����-HQ�5��
���Ta�n����b�mLwky�UR7(o�V��;�����r���j��ܘ��{���\��mGR
t� y9����~�p���ۄ����vU��w��蕮B�ݼ�ձ�7�W���,��.��.���Rq������]dĮ�A0\n�Z^v�/��#�sÿ���[+�p�U��܁�\^�AIy�E �!D�W/C����k�:h��vI2,�W�S�f��7[֠�i)�5]p����j���H���$2��z�)*6�;��}�^q�Y�5�;200U����7v������w�������X�����h�%���\3>�V���j��{}MOvu�d�2�/M1�[T�/e���L�NO�������Բ�8���Fvc�s*�Ɗ�y;���[}�j��:��6>�U�I^!� �C��m<�r��YP���>Te��3|$A�U;�~Cx����
����Á��KA"��1j�0 -�{މ�����mϤ��O�=�1�Y�������eb~�f��#�B� ?�w���'���*TF�r~I�-�s.�+��z�A�3����u,/W�����'�k�-z�"�;ԡi�e ���)�ѡ�US�t��-H2�B�r� �*��?��4U�x�h�i���bΜO��&X��m	�� v���H�yTq���^_t�'���5)�M�6��۝�B"MU�	�[�z�O#�?�@�{�`6W9������o��涊��|$�����)Yl�r�W:lu���u��Ŧ��nG6�:ӎw�-�d{[V�n�#Y"�40��ȸ�.��c��^"(��<=j_�d��=�).����a,ޫ��n�@���.T�\���&�ˠ�B�*�yTV̓�Tl�D�����wY��4�kb㋞o|��?ā~�	9�f�E��BR�&Ŕ���4z�,�26���7�����Dff'BG�صg;�BF�7dY5���A;�?����#�'���6�}��o��%�Us��i}ңɌ�v�"�\�yĊ�x.��YN n����2�U6M�d������9I�.Zf�>ri!�4��uD�3C���L�F���fL2q"t^�{��1��+��Y�&�+�;���I�wv��4T{e�F�Fb-��L;�~D;�y���-��񂊿`˺z�E���q��2뛶��ǖ�3��WD?���[l�{��v�B��+��1�ʒO��_\
պ�a�1�7x���T���^}��x�̂:��)�����'�&*�M�Ҍ_�Z�I�ʦM�Vlz0г��� jC���@��OP �4@��j&>!7�R3�ݭ��	�jd���Fy�Hh	�]�
$���E�)���$����(�_ǝf��a�
r-;������2ݚ�.��)�0�ޮ~+�i�j����&�����v��PhgVY��{�љۍ`�Mx�'dD�.1�����$(0���k���#��J�L��u��:�Mu{(i�3�b�/q!B1l!�bpF��u*/�1i��p����FT�|�+3�z���0����.����萴�aK��\���ʹ�f����$���
�w����b��+G_E9�⒠*�C1sϜFF�odۛ�������*��ʾ4~�<+%?�5��l/B��͍�*��sd�X٤F�����*�R^���$��~Kj@��qQLB�Qa���P��6y[�b�ܒf*�c�+^L���oh��ô�k����02�tdB�$ љa^ �rz�ge�~h{X���A���� ��9wM�Wʣ�`�}+��wѩ5�E�L�_���X�V#J(7t����>,��E�3k�DE��y�\+�]�y@Wd^��]Q�"|�4R�^S��D??��_=H�#A�,����i�95L���<5߬/JG�H굿�K����́Bj�`���R�h�V�X�t�kd�'�u�L*seqg�I�r#X8+]���B��&�t�ʋ��.4���& ���=�9��L�sά���a}5���H��mӴz��N,p����[���WA5ۃvYQz)��3a���C�l����f�j��ERtp��*���b�g3�w�m�4�U�OTş�rt���,}R$�?�ՍjP��4"s��j�(FWJ��7�q����~3q��(&��ɬ��J=�0Qd��;��@�F�֋����G������F�e�^_? &܇��[.����Ƭjd^b;��yֲyAQQ�m�t��i�3TE��99�s�
�v�޽x�6��ghѺ��l����ر�,�D��!91��؛��K|��jRH���N��.*��uċ�8�������z���ͮ՞�|y��� 8]	����O�Qv3��V�3���Wh����0x�3�7;;��(Ӌ�ӛ�§��b�$w�[����O���\6���=o���_�=��?Fj��j�f5\5X-9k��Y� s����{��ٚ�����k�i�w�+[�s(�Z5��T�:�W��sc{
4t�6V�bp:Ҿ�U�f2���Zs��z�G��4te����6[�w����=��-��&�)��_���-L�_iR�(0wM��s��;2���o��垿y+#�g�eU���~�I�����zF�.V��~"�㫠��WnK�`�s���n��a"��'Q]�-��Y�Ih����W�$�b�N!����<�B�����$E?�)����,E��(:��xGW�G-��@�]?�%�S�FУ+=�Cb�aBts�! ۤث5?c���*���ڊ׹��`j���҈2��QU��̣�3����26��u�z4��`���ǩ�	]�����d��и�~������SF ����������F)X��/��[qc>H8�WYO�Vh�� ��pB�;,	>af)����춀�+��Ә�p�< _���� ��NVp\t�J��*-jV�+Ԉ����]E�Fql��[���+ؠ��[[��Qm����1�p4�pU��5-_b<��	��/p��s�pu��drF�Y�z
݉�<8�4����,=��l�i8�����#����_�y�Y�B�>�?�&B�V�\�)
]���6z@��ԐeaBD� R"��M�E�����_*�q��!V�U�F��{�%��@9��m����v%#loS�6��)�<��z�Z��8N�W5�����~F������K�M�Y�"��,��]��*�8�_
�]~���=�l���Y��t�Y_�����~��5_�:�sD�� ����I%�YC���);o;�͋��UF���.�Yu�y^�݀�0My������rr�ټҿ�&���e����WX���8������̗���0�H��,���8�Y�eyB��?&&ַ���Q��;��g:��i1"=�¹�U�6��4�s�0�O�1��9ܝ^(5SoE 2�w#��5��aG�Jx�O�Y�s���<ke�&���X(�!c8�f�~����v�����~���%����V`'�ju�����E��"M�[�:��qy
o�`��x�z?/\Շ�T�\.�;[�10*ܰ���;��q�g�A���>��5\��[��H#�1l�Ntڒ��-čb�K�D��g�0�\�O���
���>5�G��Пr��j���b����@0����w׽v׭��,�K;X��`�]�tۭai��	���,����_{l�D?�)ԥ�7Z��E��s\��׬),9Z-��c$�}s��8XS�3\��"}�^ "q��Ҏ��^��m3�k�CoJ��«]L}6�Es�8�J1�X��o�a����-i�N�W֊�#`��j������^�D�z$`n��oc����K��`?�'w��p]T�2Njz��m�~��o������i����F�1���ps Ioںx;VA��7o��)��X{G�ht�t8�B���A�St����[��s�����d���$Dv��D}�_m�#]�.�Go����!�6@�k�Cر���ƥ�}�8Z=��^*� %��z�[���N�M<N�/�DN!m�1��ld�.���W5���=o�4�$�w�u{���$pV<��g뵄_�����<"�ߠ{$t~�!'�2�2���wJ�k$ ����T�#�����h����
�U9$Ι��X����W�塇J�˹��H�p��ۙ�J�[D�����[��H��#��F�w&?oC��%�L=�D�Յ�]�Y�W�=�>:\Ҁ7s�8�,}R��0��pC�m3_J���f����/_�t��,����~s�~ ?lS������:2w$��熪���Ms��r���=�t�L,ٳ��;�������'��SĔjO.|���h#ɶ���4ŐKY��~������_kn����+fv�|^�죩:V��7L�UA�ͣ(>�zČo��*4j�U�ϩ2�;�Ox�����+�UF��G~�"9�7�g����J.������He������N�~��ђ×��=���0
ar{)��s��� �H��}��J|��/��Z��W6я�[�-Rg�A��q~U�}Ɛ�֦��C͸��2f��:VR�];�����W��|�-Bn�PWy>f����)qq��B]��0w�I�G����@���_���|�f��o��s*|B��*Y"����DL�)�}�Uo�NPGO7������́����P>���v���+ٻq=[p|k���$�f��f�F4Q�m~�7�ˏ�$�Q�����6ѕ�]�$)`5�C���$tBާq^/�)�E��6�.5�{��h?T8V�c*��'�`��i�a	�U�oF��fɍ��I�!��}�/֐2�Ȅ�Th4E� �[X�,'���������.ݏ���~���Μ��(>g���惵�����y���nңE��2��0��x�!ݸ��ʧ�wG�9o����۝pl.�ڷ��z3�y~g���<-N���g������"�T��]r�h/��ۛ��@D�Y����R~Z*J�g�'����|h;�ԭ����[����V�?��?+�Y��Mc����~z4��X��w����c5?/ɹ�O�� ���g������`�]�R_.�g,$��֦�]����y�Gw���[�I�T��ɱ�{`�	��[���
�e�,{3����^_�����p:]���a��8�Rm�z*2�L�ZjP�l!�VU�˵��{�NBKS�E��1��u�>����{�ޕ�[A4Z^��/�#��{���ڠ@��fg�$q1C��S���ΦpBZ�;�;�"�iS}�����lg�[R��;} �WÎPY���_���o�:ZHܫ�����޻׌�h���&�2n����������������%}�8(�g$밿Ix<�c��� P�k�7������k@���X�R߾�W1���`[(�o��S��4u�.,IT��G9>�9��ze�8�.�@__z�y����z,wx�����0߹�б�//�-]!_v2�7T\���<��H�u9����/DG{?t��Qi����Xuѷ;L��"^��>�3��c�[k�7�@�������yqwI�.?4Ÿ�R�tu� iщ>�9�Ë�x��ym��o�|zf�d[�~r�����R����J�~sc�3�[�����H�����ް�1&��0��Q��V?p�L�g�/�Ӣ)��}��{�A�	G/j:�d� J��t�r�@��V)���eRe�ik�BtT�W��Vo��ܳ��)��(ǻ����^��t�Ӟ%JF?���!ם���Pϟ��[4I�(�w���u�o�B����}�T���납�#8yf<e��ۃ��?�n䎄n�I?�u���/Wp���&=�M�����u3���WY�;�Ye�2��l�������vS���`�ީ�E �
Z�_(_Mem��`nD�_�������%s���o(��v�\ܹ�Nu�T�9�6#ל�7��4.�ϑ5�NW��?᩽9��Zr���s(*��8D2��]x� ���� J!�^���rK��Kz/�S�� 7���A��D��e��@3TP���e�j뫥p�-�f�D��G�{�.��*�"���/_0jF�T�ֻj	2��m׌��k��a����᳞a;��*c��dg�V���$���b���ة>���d�j�2\�4����(�O�?�<k\á���
Ņ����r���#g/?�dO�1����鴍�1��E_�uɎ��*�n��<���?����%��x�&��	~A��QK�-9~��Kƌ�r��Td�/S��´��ߔ�ON���*�
�ɏY��l���I�B�& ��t��y�)�M�ۃ�;YM�����.�+�WO	��~���Ѽe1�W�(��f�,D7������=P���Yؒe���s$���/���&���O�>ı�����S��#���v��o�����~w�{����W��<�	�,?��OS�oH'\V�4aI=l�Ϩz��T���-\�&�$'�c1�y��	�]����-����۳����0av/��5w�����%�̝�>���񡴂}L�p�b��l���?��� )_��i�>��~0g8(���	��+!��}�@��^�,c��� ��l����� 	
Ɵh�T3�m���'NB�6B��z�ŀ���};���K�.[9��_�6�{}Ntncȴ��P��y�.�.K1�K�|�1� \�/Җ^��c��dt$Z��λ�381Hu��]d�<4?2c׏E� �"t�� �Q�"Yf�1i���<��6pӦWW�H"<h��o<f��ok�"����?�)Q�6��������ÿs��EC����N����f�'�s�Y\m�5o���w���WE}�۠/ /��Ms���	vÌ	�����դ
B�m����>U�o4*ȶ���fUΜ}&`2,��Cy<�[�$��}��s�J���o��6@G|гs�H�?q��&"T���Ю`�k�X�q^a���m�h�o��7�tww7J���0���%%��4�J7JwIÐ.	�FHw7�������z�m��v�'����)�q������jD7+�/3��G����g��S��;�v�����c]S-%��z�d��J��޻J�<^��n�+�:CUpph�/-���ŉ��)�?T ��$���D?T��}Y|��V���"eAh���ҽ6:^J`�ND�iӔ5��T��@T|���.�p��6�2�I�]���ʚInSfߞ��,�Lo��p/�GAk����+
��fM�� I^��̸:�K�b�e��~{A�	�'�/�*�EW��p�u�$zbg��1j����`%��4t<�`N^�.����Zd�t;Ć�ʹ��C�����!�M��e5��_���B��[�G�$�[C^	V_?�Ͱ���n}����X���[]���4��8����.��ĉ2O�K�+�=�FW.��4m�_�B�{#"����M���J�ة0θp*�����+���:ԻRFM}E��ѽ���c�4`ųK�����x�:�H!p���]����b����ƥ^$ʮjg�a75����>��{<�����cU/]y��~�������wKJpt�����̂ٹ�`X�������%r���7�&43��������1�k�"�V���&ު��}����m�s-���8?�x@���f�^�[��n�H���퐬U��~�k��u奍HǼ�thh@ǆ8�E�XԊ�%8��K8�����
"��+���J��l=1Uҏ1x?o�'�`^���z4|ƣ��P�+Xk��N��1҇=7���:��<CB��XE�!2䎕���X�4�	۲[߆v�W�_�~�ak��:H!!y�lѿ���!t"��U$��*�p���ŏ���eY��-5��HU�Z�J	ޢ�;E��1�"Aju�R��;�J������?������X��&-�F]))sƧ��X&�/U���!��& &�.����o�'ﭴ<tǊX##�#�,4�/�R�c�b	�Pp�����і��G��v�t��|)<�l�*�������:gV!��<`�@�E���)2}�_Q�Z��I'���ѱ�镋�yi���1!�PH���6J]�5a(��6:~0>�y�ʂW�wV<@Z��m�ڹ�R�SM���|���q���,]�[��Ь�ܝ����|���gdTԋ��b4j_������մ{P
㾏D!�9~���<��|:12�+���JMy�į��ط��@<��I/	Z�OͽGkh�=�Я��}P`���x���ɒ�\�/F�ҽA|����kk��i6����5
�$�'�E���W-Ȝ��L�Φ;x��D �wnn�z���_�0�:����o�W�r���\N
�w?�`8��6.�P=��>�S�Џ;q�`%�bCvp�2���Kb��
m��>:
�{�cUn�!"�dl9��,�':�v��:%�����.�	���y���W��VS�$�.����O*��d��2�&PA<��+=|;��k�tU�@���8!�����L�sN��V��g.\��;fae̜�z{Y-�C��)|�,g��鬠�kJKa�|7�Ӷ�s.M��`q�׎�|-]PA�0)�&��kb�	y�̂v� $)�ax��^�A�������䀅��a�*�GS�^u�(�匲��>�1�49�h6t���s�l(o��u��/��i�����h4L]dw����^�Q��J�~R�P̦�0<�g
>�M��hv+x�0[�ڙ��"���>܎V:���B��C����6�g��q��Ȕȵ)#���ߕ��|v2�X8;|�ߘ9O�l;���%^\*��[S��kH�&�8�T)��P7������-�o�g��~�&����.����8�"���{I�"w�Y�f��Ɔ��D�>�ϱF�a�@�\�c.a�j����8 O5z�xX�ŕ��9��3��ՠ]��Nz�R����Gg;��G�ydU��ؐC��6ېq�h��&n�pScsl����9l�웩դV��J��Y_s�5�I�E��Ĭ� $.��X� P�J~G���6���2�P�!�{%��@H��N�Zp���{��a��5S���xU�ͱ�U��F����
����j��k�q��ӵ�-3M��{��s�_Գ*�M�`^������a~�p_WcJV��gN�p9�����ǃ��a��@QW@�E}�D�����m�6��O>r���Pa���T�!��(긺Ɓm$�I�Uir�ZO�Xp�qY�ڈ��[�Q���m<� +,�����9,{t*~��lk~��T�~/��H��=!�҉�,5n��I��+1��1+�H�3�O�I���Q��a����
�c�ϯ��X �u��?_@�@��Ə�t��덙u~�Q��g-{r*���zփ�'���R�ی�pﭘ1�(�&�^���o8ae2F�����z�[R�fN��x����!�i��ڛ*���9hLTF����@i7��,���ٶ�zB���
�T�m��&��Z�F�īh��T��2R�=Ssu}��q�� ��U���D�3���S��Q/�ߜOߗ�..mxD���#_�5�^,���� ����o�c�ax!��`t�3tj��^,�nz���\(� v�`b^iLB�"�x��j`��?�I4;	�:q�|ʢ=�{��9bF5xv�>�;���9����"�����V��}}�f���F���Ԁ?.6�����=�E��c~u����O��m.4t-�l

M�b�E�G���a�`5qˣ.~���no@2����X�~8�D[OD)E�稟<O-Md���A�ހH������4�5U� �x�)��Oi��7�b��З�=	f�� �x�d\����O̥��jL��Wk��b ����Q��A9�D��+}��rX��Nz��7���4|����z�R�2�~J�a��Q�^;1V ��o�K`�.��*;'ܔ�IP���M�K�"|K}����I��н��l;��X����L/|��Wy0S��79�<y��aRR#g^��>"�w����g]d�
6����>}��x(�{�� �RF����Dq/�)ךޑ�v�Fk������9%i6���t�5���@����QPք���ߗR 8���� �ŏZ�۷��v�� �	�7�<B�m��hj�M��*׻cn ��T#K��/�1<B �f�
( i\�?C0�}dU�H�W=JV=Fš�� %:4�f�U������~6�yRR6�D�ɷ�j�(7��^F(��}�4�> :��?ʩR��?�:�ቬ`��r�\&�gB��
�	Z18�
O�)=�i�$�هj�W_�6��*�N���-��[���?���msÖ4Ҧ��F���T_�km��>Z_>D���3��F��=~��Ր�
�f��1�Ac��Y�-1�-o��;��u��2_���A�ޏ9���>�M3ræ�\�=�-��$�*U2
���i�ٴ͌�;So���$+��h��}r���e'���6�pl�¾�~�Zg�*W)-4��R(���=|�hOwV�5��/�з���P��)�������YNL>�+��Ih?/�Mz������,�]L�57r��=_ß	'��&<7��\�k��/yx=ӽम�֣Ƃ����Ӊ��,�����,��/W`��s׿|ɽt�qd��5�\0�E��q �[�?�^@�}Xyx��K�W�MM��z���y�N�ޒ�!s:K#�BH��m�}��u��j6���A�jk
)k�2J�Ko7�qE�v�Ǧ����z���w�9L�ı�]/���QZ�h�������P� ;�{���bmU�36�'����Pʂ��`0¶	��l2�CR<'���a\�@HWP��ù�40�)�| �cp�a�ҬoF�3e�/�$
W��������H�Q |���2����*�#q@�����c$)�_�̢P�gUM�uт�Z5�'��ai�>��q�}σ`�����6A���&oDG�M��#J�iF��o��m2�y�;�2��h��y�;98���{!�Ƶ�5죊���ݘ���r\��G ^��'�����d�jQ�,�WvpO�N!9�i�_:�0�r�Vn}d<�=`��'s�*���d��R'�%2e��ݺ�a9V<\�ϰ�/\����T^	+�?���l��ܦI�L٪���!��>J���(B<�A�R�S��c�+������ea������HG,�) �1e�ˁ�1TN 
���G����>y0pQF���a:B��g�1�ǳ�7�;U�]��t����rS���K�W� ]�3�}�����A��<A�ū���c):Q���A�
��o��W��\."�I,:%��/�"�C�\�tq��_t�c�	:v�:�9��R��{�}���D.�:$�
3>�_�af}TT�Ú>�>I������1z�>��;�`����[�>`���.����[���h�Y%��اM�a�U��\KF�t纙,M�k�j_)C��Z��_���F�R%moH��Ό��}YL �����F�9&�9�����q&̞��-:�)�\Rʭ�ux����*m����Sq\�pYnF����¶`�%�R�v|�C#���C�\R9ь/�Y���y�#m�[j��5�/ٱ$���e�ק`�ld[J@.P5G��M�����R4�oX�J!:��%��)(#FH�Z2t~йf<�'1S<]D�s�OQx� [Hì|[��IMP�M�Yn��Gv�"jv%��j�
,\(_9L��\������G� ^��y�x�=�r�}�<��y���j2�|�ag[�m��w>�k��g��V�!Wۇ�rXe�\�{������b�������i���oqj�
��}�1tI[ը/&K5N�G[a�𔵙��9�hFvs��ї8YQ-f����B�o��{`�z�ٍ��Q������Y�ڰUe���k�Ⱦ�|��~�n�v���N9_�GF)�O���o�~��խ�W���wBN��^[R�� �{��ԉ�zYUׂ�Ą�U	la9Z���`P�~�:�do�y���C'<~^��c~�
�� ��l�wCm-��֫@>d�*�A0�w�(���^/�$���͆�nm6p�[^�� <u��������B��|�6a���!��Vf�@?$���Rk�Bs��T���T��ZN�cO$�B�M$�������`��Ji&~��U5����&U[tu?�zb���w�ޕ�W�����5�?dO�h��sT��z��CmM`q��Pi
�%Ҧ���yaC��r�RrsA���37���CK�H:�2*|,n|��Tu6o����_��/y΁4��U�=Mh��B�b�S��ؒ�v�G�2��h�'���55
M{D��M�k� nD��?�?��^K볠[쪷�k�����Ww�C~��0=����B&���
���g��W��A�r`�i=��L-K��J�S��@��h'Y�M#P�_/�Ձ��@d=�<E2.R�
|o���{Ҽ,�`��Wn�K�Q�Ö�q}�����s�ys����c��� ������
	L�\��م[�h@�.��~ƌ�	�/	U7�%+���>���V~�DL�D�92i�Fz��4��y��U�~[��P��x�����C�+�QjC�
q������w.��/�%�{�}�K������;3b�Aƛ0�������LU�A������㭻7�sFIìK��81Whaٯ��Y�ݯ8މm9@1���0��I��ϟw�'M�cJ�I��Ǔ#��ɿF���(b�L��P{D6���?��!q�#���ѱy�g
�*)��A�~g��!-�Wv�
�*�Ty�Q[^�x%_B�4�3ή�/���-����rf32��I^L53s['���W��&�*A޽��U�&����ZK�蔘���qvd�ځ*u0|y	��f�e���z~���i��T)�,~�UK���������̿�?Q�G˃z�9K]���^�11(�d�(P
�ry�W���_!�����P�#7�����x>���ѳȱ�!^��1�9Α?'��H �vNq�{FI���}p6]}�/U�Uh��B�d��L����B��m�8��P����"1�) t�N�1�qC��BY�Ub��Z��t
�:����[�dFD�rLZ ����B�%ϥ�u|^��QT��Xl��T(�����	:�m�ݚ �J�֨�I�6���U�n��\e3X�kqu��TB�fY����*���`�.���뇇��J�)�
)[ Uqzn��S�x+�@I�=��|O1 }x��y�j�S̭�'S͟��~�u��.9y���h�6������25��FY�� �8�3c���eCS��y3sl��.|���g_]��}���`M����ᒖ��q���&#�rJ�ww���`�Q�M��~�_L<��6���;���m���ժ1}�h<O�C�YDO�G�+��������L?��j�W�鉩3��b�y���|��r�x-7�ynM�Y�1[*p^-�iл�N�� ��pٱ�t��R@mL=�d|^2ٞ�j4����s}Q\ć��@&^�+׭��h*B��'�[#��`}�l�o�7�XM�*��2���	����F�R�e�'[��CT���Gv�<���O�Mq_��x�5�ǳ�Lw�Ϙ�<s%��(��V���j5-��|>4���'$;�-ͭ��V���-R��l>���9w�,�;:����I0�PL��[�xݱQ��j�\ �������/�a���V���م#�o,m7�Y3���e�j��������hEF�<1$��%�������e��5����1u0i(Q o{�\x�}��%�E4Mj:��OJ	.��?n�=���
���R��N�z���T6��H��T~;f���l?|��a�y%�EnG��^�x|4.K+�E3p�@����"�U��)ݱ�EjgWNX)��x�ݘh�%o֗0$蛻̄�ǩ�Ə.q�[Gֻ�^���nM�%iuR/�#�ڤ��}�\qNx;$5�B�Xd��H���˥�3�(��ş.��/]-�����Tl�S����}�K�����ݭ-+�*z�5]?z8�+�0S��s�5<{r�8:U;���;,M���6�A�$�1�����후Ê�W�C$O�LZ͎��\�~��	'Ǌ���+o����]��>?@�� ʶe�Z���3���-A(2���2���ǇI��?�/-��^Ω����}���|/g�ps�SH�_-���Kr�t#��V��Z7��(H<���CL���؇��Z^��h�b6ED `����L�>���\߆��6�� 5
�+��3���4��<Nd4s��	�_���w~Ɇ�g��>Q���y�d{���DC�1_�3Q��:�mU`�s��׋�R[�������-D�������/	M)ͪO���SZ��M�֨Ԁ}5۸S��B�ן���� \q93�q1���&o48h��j�Z��"���r}��i �"�5>�VC3ꏹ4�f:N�@Zծh�O�<��)�Ȧ���M�
����������zn��+?;Oœ+�-����p�U���`G�{A��$;��E���x�J�_n+(t���*Sa��4���ڀ��|��`� oYlg�kR���z�%�����;�Q2*)(|�*!��^��">��;�}4�Վ/�=��67c|��ħ�ui���j�yd-�<Km���p���T�֖�+�kǔk�/B_�U��|v�9))X��"�~r�Dor�s�`z��o7)( _>� ��>�h��������WJ��B��r��=N"��aCMf��J���ި��Mjՙ�������vfiri��.i�oI�LE��XX6���Ԓ������馝���f��9���F��׽l+�����4=Z�<��X� �N�X�+Z[xϫ�NQ��˜�4Uf\gl���+��´ìfF�5�6��W
:�h�׍]�|]��0ÿI�e��ֽ������k^Ŕ�">ޣi�|�,��j��v��uz�2�n�?j����o��Χd^�n))p�Z���ft��!��bk��Q�݇lT�A��e����q�>ι_��*؜g}�x�1*���J�"{���;���T��H���^Iv��e���[o�̢��Y{w��f�<� �'N�r��{��1E)�rb <Ԡ����ʫ�=5�y�^&aZ�*�.��������g�&�m�1q���X�G�i��c,I�)ۗ�Fk�`��Q���q�U��ߔ�`� (3�?��Y�׶�f��nz��Oe�L���!��oݮ�;O�LQa�3�(�Z*j�U��8�����1�[��`����̾�z7m�����w���aU�C�����jOG��}1ŕ�����;�q*�5mD�$0��P��j�3�$�=c=�~o|w.�[˾�d�C!P�p��]�#^q��؀��I�VZ�4�<8�S�E�M�,gm��A���%����q\ِ��;U�}@���xk�A@{��6BN_�l)r���F�ז-4$;�o�X�3����.&��~pz��F=R�<1�>�h ��%U�jY��2;
�Έ�\�N/Q�|�����]�hH��X�43��q�Ib���*���QT���U�$]7�f����X� �(� ��?�R� t�G�'aI�T31�n�P�z�5�v��t\.�4�o�9�Y��&^�M�p}w?��ІIwUwD���8�9,'%���k�\wFk@s∜��yt���'�cc�2�W���%;�R��u��E�o�����N�z���t3�:D���ԩ�)�r]�6�/�,b��iÌ��#�HA}tZ\��m��і�1��\�X7�V��K��y�� z�Yh��\T����P����?�Y�0�+L�:����7�u&��#��yt�DUh����qqJY2���&���A\k~��q�	�РBfWA냗��K=� ���)l��/iԷ�$�-(4���<LHݪ�WҶ8&�mƔ�q%�t�m�9��6x�-X��2����z�c_:y��_]%�IP�H^� ����;[���Q���i�%Z�����e!T��S'z�be8i�k����u��A�oR�O��V5�;����1���TŢ��U�M@Sb`����
�أ��Y���8Oh)���M��oo!�d�tS��F{H�*��r�����w<6y�`��b�o���+�"�h��y��:�1CZ���m4Ҏ9���B��$A�#`1�W����I+(5���r��sO�
72�Ƴ�C#<Ӥ�7���h����֢=H���x�pU�3'�[�f������y@B(�"4x.����y3�=���q���ԄP~����0-��TZv9Y3p����}�RbcM���]�''�~L\X;��Թ1YA�H�wDP��/��P*(�Z��1t�U�u)�E�N���ai�E���`�"	��sbj]�{#��s�▗��g���"����?�3w���K������v���Y`^Q��|����4 �i�ǚ1u�%�y�����^J+���T����u�IP�ިd.�����ȫ,�Z�F�.�O�4�W��tu��7
�*���MU���_k����?(�&�g��;��H��ѽ9$�AԽ>��ݪ�8�c6S�*�A�w��2����L(��Ft�̼[��CԺ`�cNY�vo���!�3�ݕǻM��.W�;_Rhp�х�د��Z���^�(7�[B��(���9���q��R�m͹����J,j�)JP �Y헌d�8�>}	�V�m�h��ۿ�wGY>-"�~���	�`�k&�JA��{�Y���tRa�n'�f��[�����ȣ�6ck��@_��?�\��j�^C�4�&����d�9����1b�6���r�2�딶�o3�3��3�.\��/�^mH�9�5��y	#�m��ץe�6R��Q42�q<�y(;1�R�������b��	ZJ�[h�4�:�GJ-�F�Z*j<^8�N+f��tMb[��o�sX	�9p�Rǚ7繝}8���{��n1q�ǁ�iڀ�8�%S�6B1�⋆�tP������,�%�w�
�70,D-�A��x�飄\_N-�.Ւ����t�y٤ɳ�L.�/��4L�^��L��O�<����2H[�*G�%r�W���;�}�d�3��զ��)b�;���}������PBq��'�},T�/HM��~��%�<�W��e�3���	,Im��Ʊ�������~}K�������J�A'�V�Ui���#�.�i�5�f{!rʱ���5
˰���*5-�	B��r66�C�H����#�c]��n�>��+.�ih��l��s�
�Ly�?"���oq~aD8��t��x9 �Ej�C��
�eI�ߠ�>���V��uE����#-n�4��i���nB9 ��ι;<TӍ,���2���B��6Ek;nu��dg�i�5Aw�٤��N�!��l��j���0��Y�\o���k O!��Z��B�湓8��Dg�������8����Jd�\K��I����a�z@�����U���	�d��1x�P��;����zUԖ�H��S�Zvz�l{sg{��Q��x�E-HC#�o-d*�fI���e��������x#����)L�bbuE�P՚[�����&���Q�ӷh����6����d\ew��[����E� �W�,ʭv5��G��'\��W�����:w����t��D���8�ΩUUH;�m�΋D����|����[�m&:�!��C��K�.�p��l,4�s������9e��Y=�%�p0��^ňˎsp�5륬�S����b&@���+G�J�d����Z�)e;� ���J�T�����-�_*3��W= �=����
ȾJ�0d�7�+��E8��w�l�w�\�)(c�0}��\�ڋt�C�:�w�zGD�ԓ���Z�0��e/���4�bI����-�� �/h=q�<�	e>���^T�E�3�����Ne�������}AK\(ݔ������������G=5�*a?���`�g,�_��i(�~	��m6�����~�[��u�>�:U�W\�����8q?W���f3� _SCıّ�������+M`�B[��2���E�hU;�Q�.9i*��A�_fo��\8�hw-���_)&�]L�?r�K�D�&�4�P��n�m4�hC�ŉ�o%��O��c���dݧX��k�V��_H��s�����'�r�C���� P}Bp4�a�Aq����}��"NA��?��!�l�zd�;}�Bn)].�g}�iQ߹,Y�[C������0��i[�D��
�a)fM��q��P�\+q�%��-?v�RD�Ϻ��dLl��ߨ�0�-�`}B������Y��a� ��$?)aK�h<'�Wם����.^3�$Z���1C5��?�pJ��;rV����ɭ~��)���xI��1(
��8C_Y�@���A[�B�Ev�m*����-��R�MЯ�k�-/��c&�`��2�/K�9>fb	Aā�M���<��q<
?z6U�0��u�V]�NxS�k��Ų��?D95�O� ~� ��?A��7��n���O�nqrP���S�ԕ��V�<��M,O��D���G�9�#�S�R��o�G����,,#M�p#����j^6��1�V��j���f��G��`���/�0���L�)�@/m��{�.Y�B{��T����ea��N͡ٳ���[�~;�U�7H��9��Sb�lix*�ĉ��8��{�+(��6{�L ۤԁl��0j������J:����#�'H�|݂-��*�q����d#�7mv�f����sR;`Y���tTHс�+]�AG�G:MV�F�cmw�O��i[gj���.�?7�����p�!��c�D�oX�;sA�z�_�̚��粑�������	��@B�^�^؇�3v�$��š��4إ��s�sB@�<K�uB�nCW�7hOG���#���;�[y��6ņ���EfNlsw4���e�
��=F���љ��]%����V^c�� �G=!�m�-X�[,X�`W+�j������o`J���s�?(�_$��ex�ޤ�ݸ6z�)���F	l�c���4��v�q����B�����gӗ����>Q���-ԇb"1�n�t4�I����5q�h1�c?D�o����2�����w��I�u�^��tPQ��KV޲p��:�]����)(�À���j���x !Mޠ���I�E�l�Y������'���m���	���'>@�@�w���\34+pzY"�C� �җP �lqAg_�o�)p��X؟��ى�cB�;�%�_��d��ށ-�����mGY�tK�����gYx�I75�p�+��F���.��s�Ѥ���,!��|�y6�~;&Q�>(n�RXO\�|8���7C�~���ѝ�j����M<J���F���R�0<<�����y��Mۄ�2���l�t�h���<�[!�R�Жv>����I�z�%�F�˖�#�VU���U���N����f5��v�5���)��E+������V�L�ܛL�Y�у��8��7y/,N�m��YLz[��X�����y��34�'郆�J?dl�?s��6��;�w~D�}:5At<�ǙV��ӪMq짯�NE����	0�)��F	$�lȯ7�t:+ƀ��F��^ŋ4��`4�g
粎�M���1f�?@ܚW��L�����O}��#nL�D�	�KkK�і=D�|X���߰�����sհ>�w��Gy���=؋@�7�u;�.7��!)�(e��Cu�$��P0��K�j�]�
���տ]��).�ڻ��=␹ٱ��EH�=�3�7ŚLԠz�=�䀌�'��W�hF���{O��u�� ���Ã�y�-)p$z������D���v ;�ǧ�C��n�STH�_�wm|c��L����D��iy�&ـ���}/w���\�Z��5���\�[�����$�
+�J��q�j>!ҡ�Z���2k��Ҁ�>�ɧb���o?�	�RgS���AY2���� N*��,�5D�ygüN�w�bk9ɷ.�$> ���A���^�ᡠ�Z,�!��`�jh���[��B�7�SxB�J�><� E�'t�;/���6*�����`ٌ��_���ooc3��|�AU��v{x2v���
���!y���ۛ���w�~��6����x����VdTu�}�Khl�y��{��v>@���Yِ����h�:d�r�R����[�a��lY�[I���E��������u��ʹ��.� <`��a�%��!Ye���y vܲ?�`sC������_��r�QR��Ń��Y��:WI�	���yL���u�'��C��cJ&�qQ��0�ʇѲpx~p�ly !:���_7(=/�t��.p/R�r_
I^-V�N�w�����8Q>���'b>m�<��]�~�$i:É�����{mK��� �2��t�7tH��(��gq#B�"��j*ͅ汘^�N���{�<RQ߫싋��W�߭�ض��J-s�q��g��v����*O n~w�zv������Y���U�K�g��ر�~��GU��V簌@�v ��D{9�U@�X�]�`��;�e����
9?S#ߔ���sq�PR���U�@M�N���/��N��ڈ]D���f� �n��1�R�OSB6v�J�,�Y  (@�D��YQQZ	�>�CV���u#���w�n����c��B����T ԡ$�������/��&�*[��"�T�`��'�$��g'Pĵ�O��*��vN��'hjJ�ehfF�m�dMM�<tE-�T���m�z�F}-zS˛e�)n8�p��$dL鞖�T�B�DA��Z
�b�����j��5lc܅w�~:���e��8���9@៮���sLP�6Z�RZܭO��	�Y����}�s�옭M�p#1<���JT���e��q�=�qQ���^+�O����xj�ឪ?�w�rؑ}4I�z�I���U�(��͡K���\��wϛ�Z��d1M�A�A���/�s���ý �!��e2�.Ą�@�mn��2��ҷ���1l;�f��!0+��E�K��ɪ��肵z�^v/�,f�ӕ����a��S_�ૹ��hX���XR�QӶ��=Q�����4��V�ݘ��;"Э	*��Ł������S h����D��'�4NqN��ś���"��?e��H��X�B�DO?�n�r���#t~0�~|�&׍��k�u�M�=/��vz����\@�h�*U�.е��H1V�,����Ee� ��b=�"�Z��Gr�T�Χ�Y
ukukǁ�G���\� շ]�� ���w%�͕�ǫ����1�|�+�F�j`�
q�-�x�6�c�g��Fr�e���6�i}q2�Y]R}�
����U#xsM�9㻆�I��m��Wݹ��w����uœ������M��D�J�7O���U�%�H,b܀��d����kĶz��imZ�GIwO�1КC���������g{���&r�@�s����«!<H+s8J����FΗ����%\9��X$л�`*�k�� �E�G �!��T0(����o46��	�^U ����saE��$�w�g��aJ*�YA۳�������&�^;�ϫz��WFGFƮ#������1�t6\%�*�A:���$ʥ�6o���Xa]K=%/r?!; �ϗCx�H���������f��/i��i�Gƣ�W�Q_��I��͙���4��"��e�:[���"��"7��I�� �$�����wP�`���_T��"�6"fo/њ�|����}(�N5�Y�Y�%��"�w��L��~����Ħ���S3���u�h��n��x�
:87���<�|��:�b��v���oD�_����$����[g������B��Rg�&��և ��&F;kh��DZ����(5(�_f��������dZ��'�����u�WVִ�,����h	�l�?�ex��n�g��@v����+���
g� ��ED����^\0yC۪���6�aB����uFi��ޒt��B�k�4+j[����ZRTq1w���'�XK�i����i��+.�=��qW�r�BU��ы~[��U����'��iVi-SSGd-*�[g4��H����7���z�o����IW/�UO���=��[/,�Tƿ#E���l��%�/�Ԋ�O���?�~2S�/U���z�i�)\g�w��=3��&�ɰL����{l�܃�яƕ��CO9#ÍL�j�#�<�E1�t���-���+mI>.���\�dT�>�:�4#��"�;�߰���Ӽh�QQ��r��t���q��k�c�W]�����3��Q�^���t�{Y�]Аf(y|KH7���k)$2��W<�.���V>*���3�d��<��P�Ȕ�c\�ǀrQ��S�����w����.#LѦ�}˰�)��D�o�&�ٔ���S\�%����{:��D�s�Y^Xo��C|09��ZP�<l�z���^�Q��	V���F��'�PxT�����n�m{X;�]�4e����+(K� �R:�}(Iz�\���U�-8�Y��X�&�r��[�P* K��iN�+�[pT?E׸��5��DЭ���y�e�MH:��x-�l�49������0�X1.�e��#�ܶM� ���a��O��h}��~cd��	M�����.+��0����ۀ��.�7�&�4�e�"�� � �����DC�F*}��z�>�]��NNW�Վ�-1}�����v+�_m���-�5��a�b��C�34��?�.�{�C����6[T�8���:#�)�-˯��:������sM���ڈ�5o)���(o�R;m�	���s{x�7ۈ��zM�[�^��zW�����(�b/V6�%�V�r�AW/�9ɑ�}�<���7��T�cƊ���^���	2���-����x*r�yW��U����ϯEU�	�c����n�-�b��Fg8����'	�	]������p$ƴ=NxKo!��E/0贤�)_�B�߆�������x%���<�T�u3���ls�/PQP�3��@$}k(F3���"��v֬��<����;��*���@K�|�տ��B�Hb���5z��:~#c���KY()Î���oTs,I30����r�z�������A�Y�5��02��$ޅ!�ش��Fd�����P���a'�5d��H�����w_��DnxȖ�3 \�����{}}�[ru5۷�u?�؈�M(���39�2=M��#_7��r �����b�w�ɘ<RV���Q�35j_�����S|��s	.��eIڼ�����k��E������}�̈i�пn���Vc��e�����ޜ�wޒ"��l[<j@�L~�W"ZT��F����2��l����
c�C���x$㪟؏Q���f��+Yȍm��/Rpv�%5�7�����n��!k}���o�[�U���3��m�N�J�]@A��������Х�=� UDDz��Z�" R��H��Cޜ{���;�sތ����מk�_Ys����{3�������Yn�hF�?�m	$+�O�
X5t�)�q�|�#3sf�^�ǩVxl�~�-�����Pk��+�Ǻ��^q�O��:�U�I���2���.�ܙ�����?#��p��5%�؝�{��Qg/�h��s'��<��ʊ���ҒO0y���n��$��)��AF��3��S��9X^�%o�	78Ow���3��5�W���&�!޴��iki^�]�YJn۪������]AD$@N��|7c�.Ѧ�_/dӐvV
Y_�Q����M����W������C��T]M�-��0��y.G	!˜Qj�v!3��o�N/}VUş�ȏ��I������PK+vO�Ⱦ��De-�~?�~}���L@V�����f���=?�J>���Œ"�}tՖ�'�áR7��kᇢ�R(;b��7�3܄���?~������t�8l��R5�Z��Z=m8�F�O�OS�E���ѮC�?Yˮ��އZ��b�"o��%�_�W��Ҿ~��U�}[�������sss��4���*�)�3��nO��Rj�cz7��b�b��F@Qs�?���v��Q	
�m�l^�����ؾ^ˌ����	Ȳ���Ѩ��v0-À'R���1��Ϛgy�ZX�T#H:�1`��y�jL��Sc��M,ֈ�?k�4�C=�OZ��wI���lO��DBw"�mM!{���/rj��%�!^��p��YK��	r��?�@@����x"�P�M폨ɯ�g)@��R�������A��@|y�~�L����+y+ÜK�ڍnw���Y�;���\����C�R}���=]���u��w�mHo�g�\:<���H(B
�#Lݍ�Q�x�^��<�w��ف����I�!e�����%��������.�%B��H%�8�$?��-$��u��z]DH绿~�16�uB\��#Dzc�|0>�*��+�_*Eӽ�??����c����V�z׹�����cNy���Q��o�c$���/�
�9^���^M���&\2��%��z6.��4D����a����^
���z���*����W��	II���|�z�	���|˟�&�g��a5@r6HS��e��O�=!��i���[�d��c�l�1��\jwv}�S=<U�zV��]�HE���ߡ)��rJ~{q����Qȁ���Y�"�ܧ�ew��a/�f��Z�LZ M�ԡv�����D#(*:�S��׎'l\
G�R-}]�#�C�Ici�"vn���ٜ��KzzQW
�1�qY}��0���Rp>A��c`uſp'�ܫE�]%�dS�to�@��CyQٴ!��w��C˴��]Ln,b�zͱ�Ed�R����m-�6BP����5* �h_�j�Y��݀���R�?��+*Z����%l�(3�b�0��g�4��'f�Q��?^�\���
��K�~����@^�׋:���,�����/6hH������O~?<mV+z���_�\�O>|k��>���O��&�HV=�-������Z����2ܹ@n��A���_1���_ۮ"|��5�Z�ٍ��Tl?�ݚK��<Zy��=ە�y��O��ӷ���ΰ6*i���T�8�Fc��rW�9��ޝ}(��,�{lS�k��g`�����ْα�}�~�Z�ia�w�5���@<%W|�1{v&&��`Q�&ꥅH�F�h|��B�(�O�����p ���y��WԹ
��d��K�$�3��	|��L{�)����ک�k_Y�)�Mɓ�TfiJ`A��� e�T��o!w%�JARRz�FAo���c`�!�d�N�S �4��3��<^
f8��E�0���X���Knßʠu+���p���)/�w�x0�W��m�~q����T��6���a�L��46��Q��V��/�`~Я�	��ʶL�~H<h����[���m�NN?�밓�D�P]lp��
�+�B��K��$~���~�%A=�S���L���DP�*��� SF�<6c�����/�Ӝ�I����Z�%ͱ_�A� �K�����A�5(4��p��;*�g�������V�S�Ve�淮ݐ��?<A�<S��� f�7\t�v,��?���� ��l\�%/�$��fFhk/`W�*�@�!
a�i(��+��=N�[�]��#k��t�F���}�&S<�������*���_N��fP�z5E�Q�z=�S.M!���s��(����O,X���H�kk�������O�0�xPr0�d�"�zCf)�6�����	v.�&�z����`���yST��d�y�I?��g*#��9��3�nC�Ⓚ�9t3U!^觵NC��v��ݽ5Ͽh�f�-����0��/<��W��D�>s���3��<M��d���33����k<f�-��^��4���P4�z:rc{��2uc*h�)�B<0���U�EjZ�oUF�?�`���6�`�����:�=����n�_$������
ѽ��^X~0��BA7q���sj7�ž�9���u�J>0�V���G ��a���F�⽚�U���ԣnv,J�r>�GQ��E!n�.��x�:6�<���	����'o[���<X���Z�m�z�8����J�]�tOGW>��)L�Tos��޿E��h��*�xЪ��>��jՆl�ȣ�	�D���>6�ևq��|>S�Yۍ_STAG?�U��|j!v�P6]�Jf�u�K^���hڡ��D�?�rzB�,���Yj��!��d���ں��wӹ@�Q��}���D�{nk�D�c2�4a�U���,T��ۅ����9��B��S�gZ�)��b�X�߈^WAw܅�HI0 Z5�cܯ��&9�%���%�ވɑ�j���{JTUss�ۋm��ȿ-�w�ޅ�m�f��O2��J�3��i`	u�;�[�$�(W��U�^}Y����A���[��v��fdh�hE3zO)! hl��	��Ⱥjj�z�5���ϮM�q�e���Ҹmq0`�j@_�����N������^�/g�Ǘw`�ӯH]��Ynu7��mu��P�սMD&ǞO���2�h��ӗ�&3������#��5��-��C��Q�8y�j���z��4�t�q7%E���aTT7�����5�L7�l1����,4���XU�
t�~�e
����mS�to����U�U R(p�]V�.�\��}j���k�@)X�����	+��GH��Z��ж��%m�Gu���j���-`9���.z0:ؤ�V�t�C�٪klIG�����, �ti�T���&�U�=$a��Y��"~n[y�2V;�6�@�_�Bb�e�;��ĺ|#��A��'�[>(nl���$f�ϊ�ZjK^~�R��wK^�#���Y�7��R�>��|�����[<*%b{����2���e̝*�#� c�xo)Y�z�y�3��#���U��Y��g�{R9ԧg���U�$�#\�П0}����Y��L]݉s$�s�Ϗy�w�/.g��m�^Py[m�W�G�I�c��)��Ծ�[֗��Q��,`hOL��t�rh��؛�R.}^@@���h�q�!]#�:Ҙ8�Y3�欺 q~��ALs�t�d�%��G���`�ب�]���r�yD��($�.�P����V�!��*��3 ��a�<��w�\
�i���ȯ�'�݄�ת_�v,q����ݟ��/����?�	y����ǐ!H�N
��&é��In�yD<쾖��U���p����E����C�B�H(2���45�)6ӏgބ�Ù�	����(K��^���HC|��{�zV�L|�=��u���С�:���l�����֥�blf%�]����y�>�;z-HGM��I�����bq�i�`�l���͒��*�Uh�n��ړ�wX�p��zW;�H`/�h��Rt{H´-���z�GTOc�t^�Zhp���;��S1\������b��,��t�>x��-q%�RX��͚�X�q��t�Ÿ"�0�j|M����_�`r�x�EӉ���C=����^G0O�,ȧz��/��)H��fT�<u��7�{]GŤQq�|�'��e����\�&(�A�(����?�A�Bw�L�4w���Z4p�Q6�������^�@��;j���p��/�6���t����j��,{�����n�Uy/ȫ,�����_��h=g�P�ElW�"1����?7592R�,a˒�?fP��`�ՆG0��o*=��X���j�({�Jv^����+t�\��~��S�sn�]���Z���������dI09�5j�:l��y�x��/���7<��r|�Z�[���Н+�Jv�b�Q������>�Hr�x�o�G�Ϟ,�=���/a G�M�v��9o�D�;X�(i��|<alP��Iqt[E�<fk���DtJEGo�6𐔇��P�Z&�C�m��e�2�]��a�T\�E�j�S3�������;��N�����2�,a�S��9�'��4�����u�S��;"I��MM�!;�!�V�N�dҵ���$w��B�*�U׌�c�'���4�l��2�)��_V����}K��M�����i,�]=g�F)`ttc�i�5$z���'/�����L�\˔'���c�V\��KjO
���B�$W>�M�9��pY���=tR���k]�g�_YH&�ˠ'�Z���)t%O�u>��tƓ�-��eծ;�	��qo�\~��)�����S��}
 )��
�]\�k]�=��`�g
�qe�������B�Z��Rps��~�ƻ�����,�K�;�M��#�M�(P�#t�h�	�:�ۡ����3�M,�팂�$�� \ct2��+�'�t�Jj}��݄�|S�>��^e�+=�rJZ[��ZG��3����9�$	9���a$��4M�iF�������<��{�?EM��ۈ����������uA�"�D�#�t����Q��*TS8��@�$sjr��d�*��Lx`o7�����1;N.��L4eN���ͣy!D�n�+�jH���6/Z*}��w��}˦&�I,vH�����_�h�*3�;	��S���M���,��z/7�5jM��(;2��d?�"ٟq�t;B����j}ADN�-��X�ɎY�����v5Zg���͓��"2�5�Պ���u>*���'�U��Ø#`���n��������
F쉛HrS�!I�%I���ҽ��C�`Te���K��(F0$�*�5��>q�,v8�h�:������2]DZ���!U��$o�΂p�qV]4���=E�.E	��&��3l��
:o�Ǉ8�l��pO�$9��} �ǀ%�Ɏ]�&8�j�ɐ���i���O�o�S����mc��)h�
)�UX��`�7�<7)-Kr�㜰��lqM�o��غ�䠲�̋�^���{���;����U��:�}��,K<�F��:���K����n^E]<i�v�L�S|�0��^�Q��Q�k��k����K���~~�o~����xv�ѷ�4}�[��M�$HWaSQ?����쵇��8ƹlGV8�Ծ�u�K�v��sY��%$|{s�Z@w�4=� vvx��>��}<�
Q�F[9�����?<��ڲ૮u���:��s[�y�*B9h��3�#Iv%��\C><)r����?ug�aу(�g0��O���8���Jz]���@����c%�&pj������p�<��&��U���z����� �;Ln�<��T�#��
HFKF�
en�����@ۉ[�^59O��]��q����_^�4�@)Bza��<��VR�^~��K���7���Lc�vf����Nl%x�qvX�90 Mdo%���r������1:l_o�m�*\Tu�ͫk��8*A�l�C��I[K���{I�j��"A1��%���Z��P�����O򙡼�l����+�X���p�	��CO�,(��"4H��q�=��!d��1K^bT�Q݀�U�Ȯ��eN�Ý��B���7�7W�t)�$Y��4���s���G����s����f�=��k?���=��M���q�n%X`8�<���F�Eh`.���P!6���8��"��2��^_�I��9z�,M��0,�t���� �9�	(m]��[7�)�� {a�̨.�dʽ"��hu�	=��`��#��?�����,�^��C_�O�V��?1�-CNڀ����J!���;+�ɷu)��������#��D�/�ﴦ\7�n1�G�q�H}��s����>���*�(�ŰpK�#��ؽ��F�pur��e�G]A���)��~�]�Ŝ���R?T\U���a����9a���
U���%.���m��:��#�^�'f
`yϘ(��>p�?�'k�H���t���	���A��pz�9LA�!S�[��+)_\^=+2iQ�d�.u��p�T�&�Ö��"��Sr^U�huU��%J��n�*�~f�F�=�1�>,ݗ����|nP|%�����t���g�H��PX	z�X=�	�B
�|R� iYq��q��խ�!r\���*Á�bpf���DF�������2MXtx��B������Zo�/<��e�|�(���kS��D�;��z�O�����s��c�����t[�g\#�����=��� =b�
��0g�u6�(���"��v���9�'���f�='���@s�-��b7�W�샍7�əcW�UT�m�^�����K�8�Z@�$�i��yԅ����7J&��0;�	k�������pݭɪl;�~z����2�W�m��hbR�L�a5�2ﭖ��d�̼:�P]�mQW>I�}�c�C�A��p�L�+�v��W$#*l/0���"%q�	R�y���3b��������z����_��A-��[�A͈����K�yq��)墳9Q_V����i��P�)&Ś��:��Ŋ���ߟ�N�[u���t���-;!u�
2f@��	j�sbW���wp��=ǆǺ#�qŰ�i]�hdH��l��t5�ˏsܰ�N���\�cq@nǐw�Q���hS��1���-�(��(�s����lʇ��5�r�/�ʦD���R�2R?Ej�(�P��s�VM�B�{��E�ߍ�d��)[��l� ��{� c���žϞ1Q˓���7���h�>n\�,�QOzF��VW=d�o�Eo�M�5�Np�D�Տ�;��5�S����j�6��l} x��E������=�B���j@M��҇�C��n�<j��l4��]���k�#C�<��m��h�ŜWX'
[TU���J"af^W�W0�ڬQTȏ4̱fyQ�c�HH4�e�O��A��F� ��4O� ��q�1���s���_X":I��0�ȳ:Ǖ���L����wV��Co$+Oi^��۬>_Κ��@��B�&v\qij��׹���΂ۚ=�1��ˎ��xY�c�ZL�el�z�!=H#�SA9��ƌ��#0+g�{^������@�����aU����Gf+���%��R�ed�
)r]��R2�2խ1ЁEKZ1�ց����t':�Қ|#�nf�c#�O!(5�`X��R���6�1b�rU[ǧ��]�V�:���ѫ3�Z>����!���x	��=]�R�l.�%���]�I?��V����
�\=j�1�}� 4���g�*�{j%��C��D0�<�ôػڣx��WQv����0�`�[W��
�C�Q)XL8n��HLe#~��� ��v`�U�����&ސ��bn2EJ�B������,Ѳ�b�~�x�)o-
�ɖ��&�c�W�PI:�f��O�V�����+1���A&$��;L4����,Vl�����Т��l� i��&�_���l[����zV�����|d�o,���/n��c�"�[�Cp���l�de͜�2�ǆt���~�朓�횄rGԂŁ��F�j���ٺΉ�n������_�YY�r�뼨 ���.��o�G<�R>����d����1�L�?w8f�PF·yr��q��B�����up�B^�aB���P��7�1��2�55�G�ᘋ���e�,�Z�Y�--���bM�ˉ0�U
@Ep�tF!�s���ĩ�r��_;*�ӂ{?Q ILyEĸ�nZ�K@�] I����ϛ��!����i��R�B.Q��k�w�l�k�V�O��`�����,�/��N�db� �������t����I/���s����K"b��6E����u6�D�yR�
�C����˺��7u�&]����퍃=z��uEt,���kG-c],� 9yG ��}V����FԈ�oR����b�+o�`�i4�����Q�:+�4�E��7d=���Am{�{!������rAý�*�sl�5����w�d�j�ݪ�<A�i���RK[�t�p4��N��*Z�Dy�Ib#Co���p�ą�o��Z����hl6�-�F��s~��{��>e�ķ����OF,Q������~�$C�u {Et������*�ăV���y/u�|~�ǋ��,�m��!)"��jiÃ��([�������0YDA���垅f䛎�Ob=��5��ا��qy5-����y��p/�e�7�n	S�9ֹw�)X7
d���ޣlz��{9��w���=MJ��5_f�������0{��_���O�pp���"�F=mlMa/�
�<i�9��g��)O�n��Ǿf�H�xd���&@���qۤG��~+�q�u���"���rQG�(��5�E!�Q��`?~�~��
1Q�H�n��Rm�s����$�$���i�\��Y'i��4�(����z����p���X�bN@Vp��v/�f镌C�.3�"�T�um��$�p0��~�o�7,�K���9Ώ=�VL�|t6�8K$+���/f{���fuX�ך���J��͈�<a�u�� ��]�B���ƻ&dx#	��߇�JI��s��W�)f�H";e����Ŋ�{�5�m������.$ Ğ$,r&�(�g�J���]�߭���7"�O?Q�O�R�"��=NS���0��+ p�J{��Jd��m�X�>��=zߨ�����[ ���*ח[ oE�l������rK������W׀F�\�A�3����f�"��^]��VT�vП���t���N>�5��rFZ����Z�M�[�~�>����:�h6���'�D�ß��?)R �h�|]��G��}eîHW�����f�N&�VC}���M~��s/[>9Z�G�a?��2oÇ=�&ں5�gX�F�Sg�i��[�R� ���mҮ�e���]4"�Y,I�%������
⊩��Qt�>�����$������(Ģ����R�z�Յg�q0n�Z�ĊE|�K�DN�,�M�O�U��]^����&�V�}�6A��Vu_Z����7�`�u�������p`MƯ]�M�K�wr"�7��χ�^�W���A
s=ͧn�r�W� �OY�%������ٌ��|�jْ�W�˾ �J:�����z��f_���hG;^?S��9P�����su�TI/��n����^��tu��{�)Ư��躻�$��Q����+M}�ƨ���|��M�o�;J��E�On���Djd\��I�$��s1�Y3_����Ǿ��t���H�=J�ܚ�7�#��C�Qb#X����b� �y����)�ˀtr� Aj��[��
E�/P��ruf `��K.�74��CX�T���'�[f��ז>?r�TC%�u]��ub��zJa�Z:	�X�ӑ����� �v��+��h��u۬|�>~�f�E[���ӿN��jIƺ���s|��n�t�X��hxJ!2R�$�M��5܋�*e��Rms������jf�K4-����`"���\�A�Y+|�����#a�/?"�X�n���ƅS���[�Tw�H�	;Y�i���1$��V���g^Ȭ���@��2��1zRv�����@�Zq�]m�6P7g���,.���",rMlr�D�s%��!D�2�P>��ûT$���P���p[(u�v(�m �l�Xy�����	��_<���N��f@��,�eE�޶4}��Ud��o��V�ȅѻV (~
5γ-`��a��,��d�˸�eZ��NAR>{6(]m69�je���n�e&�$�FU�w��)	;7X!^Zz����Ic��y��dͨy�^���|�?�6ٜʢh�F�0�ԆEf&nm^Y!mx�#��Yo��~^�#����7�E���$RBfFP��;Kri��(�l�^�G/��Ӆw�������F�f�38H�atA�p"����|��3�}49�E�$�R"0D�S��c���(�?sZLdT����ٛ<���0g��k��p� �����ry�'�{�ʷc0����y=�h������0����l�.��.w�����Xc�yK�O��~�_����Q�� ��+?���.8�voJ/�eR4����qP���gYTt�,��4,ޏ�7B�Ks��|���ih5�G��M�ƻU)��

��"�x���k:8��m�!�H؉eH��'�oW"h�!�s����d���,�q����%���2z�0�g�m]Z�v'.��H*0�IR���aV?��IE��xo��'!�0&�U�ߨ�<��#�u^os��M�=�ߣdr���il%:����>c��|
i��n���_r�|���@�.JJ��?��_k�N���KH�>j� ُS"��צ��im����ib��tR�.z��F,Ȉ�\�G�]4�ai�3��<Rڠ��%�X���\�_���3�&��A҃!���<��rB��z0�I�J�;��E���8�)�ƺ�0����	C���7����E�a��n�C;�"B��#������$7˓ͧ�~Y��_?7����ҧ�MîV�p��,�q���Ʈ�)������0�N����[���yO�N�q�=0+*��I�T2F~�!i}��&)G��_�$�G'�j�Ξ�v_]�H�b��������(��I�Jt��b�@S�bj�Ow����:D�Rz���C�;H.�+�K��ۄ�
��3��e�� QL'0��o��H�cc{q��o�^����xI����{|�vvE�q|>�B�m=_]:���GN�������!L�0Y�βmt��oT{�Z���m=F���w5?d:y�j�Vۆ_�B��aK���
�s{�R�d�-��΍��3`PXiR�(�^^୔2*W�YD�彛Y7Z�0�Zߪ<W^��6��C����Nn�W��\IWo��#-5p\�_ڥ7Ɇ�H%����pϤ	��k:�k ڌ��凍Ig�*�E�b�Ut'\���<}w�NڐN�H���O��̼�4���t ����g�<�����nr�c�c*c+E~�<���#PժgA���TC�Ũ,�h��&}%=�������B��K=zws��8�q&��#�L�pU��q��	d��]�-�ѹ�9YXvp�㒣k�R�M�;��4�fsT�h���4��N�v��OVgA��&$=c�Zh�����'i�����WD��b�h�"�'��i-���"7_a������,\�����t3�
�u,�O���ki��ɥ�}`���5e6�~3!��OI����u�uѪYWo�3���H��:r]].�40J�bn�Y��������;���`f̱������0�����J�}�]�l��Q�������$�)�cA�8��(��y��M�[�_A����#E�*�ϛb�GWd��m$������"�Vy%6O�9OB��$�w�Pe�G��ܧ�	7�d�>�ݼi���z���%����d��2JA2ǩ'��P��K�(���9�xb�j��=�WUk�V��2&Y|+�C&�煵�ƈk{�)]��"��M"cdiUS([�z;z$��P�������r4�`��QXK�W�_4�p�WV|�p�)���0��#�<���>��\
����h�#I1&t�C��-�k�0�mi̚��q�M>8�V��f���[D�����o;'�����Z�[ANh3���{}X���҃��{y)ӽ��gW�,�DɎ� �EES�{�tz����	����2.��F�B���A��z�=
�]J�Ei;	:Eْ��˙�pn�U����|�k�T06���'ߓ2��L�8	��[鲋��sQ =�%Rڡx6��r����zQ�|����uԺ�W���Ò��ϙ\�P��S���"�M�=�{�d�$���m��R�$l����H�ۓF��n��BN�E�,y/�N����Õdb�9�Gfh��g		��,#q��HL5T�r��T%mF)�j��Y�.����]խW�gՕ&���8�����*#c�Z1��ϮKG�zC��B��������>���˸��j������,�5r|c�]ep�5�;�+���Օ�V����F ��X�/����'����wV�����K��*��V�5�ļ�˪�8�G<u�/$):�8b�ܑ^x����֫heѮE��恔Z�_�
 �����p��A�>�C����/������PX��S�,�1k��LW�:�����pK���R���ΟƅJ�@��W�ϾPb䥨�H�TD��[A!Tf��$�H�W���()��ou!����ܿ�b����������|t�3Y�[��S���^�0�W��J��g�F�����D��T��x�,lt7��l^]s�͊�^�^��ݞ�u+���4����I"�d`�Ԧ�5��w<INQE�(���߀�H�� ]W����$���6kC����S���ֹ_��B~CE%+��h&�y�Q�p�Y�Ӭ��&ܦ)'��[���q[�/R80A��Lp�j���'uϙ�f�ݞT(k��r?
�
W�~y�*w:�������}�����Ãդ�g'E�++���HH�}���(1ZZ�)�3>��Ƣ������旬`Ӹ.�YY�cmM���ڮ`�n��0I�C�����Ďh�^j��E�BM��:Пn�J{�`�Y°��\��:� #��1�w���>��-��5oR�6�Q�|��wx�!����$$4uS��U�:���8{�@⪙>�%kֹ8�m����[����,�G�X㺐II�TCX�KVhT�E��#*SM;�\�������CAz��ɌR�[��L�H3��qS�:��Mr]Ӱ��^{���mys�6ӕ�^߶(y%�i5���~��~b�]�����G�c#�Ý�4}��ՠ
��5'��(����(�[!��PCyϘ}3X��~���N��{o����P����џ�.��v���I��z!��9(]y%9+�'{�*���[�'[�����1��f�-`uz"�?�
��^-J1���t��z���E�����bl�h�k�s�^v�5��.^�,'4��ӢK�֥�	lp���0��7��+����Iӎ���H9c0!�u��&W�0p�=:����s���0���+s���L�U�l��ɌV�4lz<������-HBH���
Vm�S�q��O��˶j^������.?>��%�i\��Q���m���7�m�#\%Q��S(�q�;���J�D�����A?$A��U�^�(�T)�{��蠼aa"���)�A!@3ըY�z�I�������J�\:�󣴷������~#��}�-�\�7��A�M��	����-����ϰoQ�φN"	�������=z� 6T.��ē�v���Lz�j��v�x����MyS !��K+�>�Z.u_�C&�'L������K�$�g(��_�Ԁ�!4���J�YV#m�M"��A\b��D��_nS�l��пJz	��2��\���ؕ�;�������p�Q�c;i$�� ����b���b��#�q�`�Ja�:�'�|�[�r�WN�,	f?��b��Pf\�t�l?����%��Λ��Y[&N�|��_ԕfOD+q6�-��c��_�3�:�3�>�l)7��;@��2�E��~�В��s������x�wp�2�w�Sl�BK�e6�^y����޻��h�/E�!�	�_ N�x�g�R��(��	Fȉ/��n�^�6E7
���/���T��e���������|Q�d~��PCC���aC������uΒξ	�����@"����}�{}=�`��ͽ��|��w꡷p�O�6M�r��-'w�ՍH�c�@	�O�
��Ƚ�5��������M�7�v�>n���V{͌l���9�,�}!	�u��
Z��6Bu��6��35���h�fx�<���:����7��
�&��
4Ƒ�?�nߏ^� Vd��{6>ķh6�l��o�5����>f��2!P�5V�>p�H�U���؏kBEQ�x���\TsQR�����Jla�/7�/%�����¢��OU�n/_�������|{�T�iA&R�$����{C�Ԭ;8 &���s�e�u��x$1�ʺL��!V�3\8�B)$���~�����R�GvO_"�^�ӆh�	��P�>+��F=�y��';!a���o�	����8�"�u��ߔ���(�2�Z5�PK+�X���b�X���7A���.�T���u��gԭ���~���˜2#��q'��zD2��#޹�N-�0^ �]U����o�/����B0J<�e�V�Zqm�^TC�G��բ��o)�9�@L}�|9����J5�^�V%�!3�����5�c�\��2����P�^r��}|��	p^����(}vD�bkYV�B؊@�'PQ��y�
>�[D��ӵ���ܔ/:��^)�|pc��S�q��Di�s�f�$����.�3�o06z�e�cm�<���_�a�;�i�Uɱ@�qK��P�Zl��5�=���ĻEny�;�N�OvA�Gvk�S�ѥ�d�/L�P�Q9q��$� ->������N�~)����?�P�AFl��f��M,/��{��8E+�L�K����#��zKSy}��jQ�l��hj�[�e_�kJ-K?�|��e���}.e�����B��J#�G����(ͽ����D�B7���M�����/��l���eR���9����Q)lk�B`E���n�%@�%���|�(���{�/��� M�()�Qw�3���315��
c����b,�'n�e�eJ���[��������?K��`�4���v
	01k}ы��@ؘ��F������Gc&�w��Om����<8�U���ɇ�䤤6ǏjMġ�:�����+P�Ȉ�;�$46l��~�+{�%MA�,�rA-�vV~%_�����.%s��іMk���{��6]�B���_>��]5�w�u�"%�S�GQGk�Df�s�-��<���H�u��ʇ��7� ����ե��I�I��?n�i�',�'�ay���V�d<���%���L���
t�$#!�]Z����[�b�Ԙ)Aq�/�/��-���~��[�c癯�~H���XK�֫��߬&IQf����,P��ߴ��τ2Q
S'��=�|�ä���=�(Y��]�Y��/��.���(�����*ϫkMS��B4�3٦ق����D]�Z��B�T�oNM�N�;��W�����/�'��i��,�g��.	�0!���>b�|:o^������D7���8ZbW�_l��;�D\:wN݉�URG��yxYT�Ļ�$�#$b�G�OZ7��Q/���٦�&���E���?<�;��ļ/�^�^�����N��'�/Yvh���g���<�&AYwo�ji�<�O���K�E��K�NH[пz�1��3�����Q��z���F4/n�V?)!B8
���6�+���N `]��|��f���p]�c�(Fv�T~��~�+|���#ׅ��R�U���
�U�_�{�r��r���)1`����&o\)�Lbv_�F�k>,��eD���L��q^�U ԩzz�1sk�7���������Y�!"ځ�_j��i�r𫞘�ʼ9���׿�bB뇵�Z A1&[t>���x����j�T%W������R��-�z�Y~��m��%��Z �/y�����˅����;r����]����u�Jv_�㖎![mf��Yh�A9u�Ph"�ٸ�ƽy?ɓ�\>$`M�a�:(�\(3�	;&ro�.�!z�'��ޖz�+3k�����r�|`X�U�]�l1SJ|J�7]��r��,J����r��f����A�O�@�/t*�o�:x�pM��G�v�S yrQ��%]�x����J�r����_��kwLh�� ,ֳәm%��s�&@�0Lp��-��}�iNx]|8�ۨ�$1�?��3�w��������/��W>�<$�X0I�20�ǃ���>͋.������,P���A�Q%�s9����vq�UKe;��J�`7��-��f(��I1#Oxj�M�s՞����
����E7{ '�@,s�/��ǂw0]Q�B�^�f�m;$�Vno\[#-Œ��gڠ* U��}">��6�����nf����M����&��9���K���55V6qEq ~����F�_Z@X�Q����m_��%��52��ʧ��ޛ�wh����s� Fb	��3��8T�>LU���ĀQ���B��� �n���:�������V�{����fۿ[��m��ԪU��^�֦���v��&�U]F�-�fQb�إj6�$B��4b�q?w��s?��^���:�����<?�X0���Hc���]�;�D���6�7��R�Ne�^X(�܍L�J �?>9��$�\��B�$US��M�&�
��@�f���g���].��:)n�Ǒ�."�i�?6�t#��v������
"�S��[y^��\x$Df���u�-O�	i�=���G����0;��k\EÑk���/��*��8H	��T��[��@Ff��-衫
M:��+���wض�/�z��_yH_&R�b��+N����P���n�R�_�[!7���d�:�";+]k�'9�^Q\�l[�}WA�ڟ��u�K��$j��WMCг������I,����|�*��`"��Bnk�����7��Ui7Ēnf���o�p�k��I��H�H��2�l�MI��n�^b��������r�,�.���ĢY�ϐ�k���Բ��G��7ן=��o ����5nm��i�t�QU���[�F&ۼ�}��駷]�l�݁�]h�3�DכeS�VE8��\0�&7���gYE��	�,�Q+�~��_�����L��#3_|e4�f��`h&���_�D�K��m�Hw�=�#}}y�ddO�ֺ�t�_4
����.��N�zB�!H��s9��Om$�6�j�Ch��&|�\��c?�b�3`o	�6;��O{�#"�^ڠ���ң��fV����(��)�v��]�Hh@�7��]�\��H�;�D�0��6�up�J{G�Sו��j78�\�B~dvGL�.82��]�(eHuA�H�lyF%�V'�o���%��;�<�����͒�}���#�1�o�f]� g{�@n� (���T_���}�alg
)��"ªLD�/�l��iM��xa�o�-�����"�yŗ2�� V�%A�\�T�~S�������������Σ;>k#����*�喡��褿����Oz2K��z��qj^t�&{Q����dp�i�G�)�
87��������=8�N���!3[��%� �����x��|�<o��E�m�e�~w��M�,��T2�	up����]��CxTl*	r�y�C2�kŽ$K&=��-}C�}�*��0�D&�[T�Q*:;��sk ��]YbW��+2�{�<Mu��^n��(I��R�	�禦���:�x��Ϛ�6��)����>��Iw�AN"�����Г��;�G�i�j�00�˥��q�R�6#SC�ǅFf�<�4,I��8�_@4mf�pNDTq}E=�~�n�[Ƽ��cb��1%<��ς���XB6Ǆz;EɃ����B���G�����>�z2��H�өL�Z���/˕�4��<�2���#�4͢l��
�T47�Ec������w�������W��V;�O�?��L�=��`1�'�.�t2�63��=��>ցf. g��x��,*���va>��ޣ�kY�O���_,^�M�z�c���e�#�����F!d�$�n ^"��ڶ��\hC���I\Y�m�'�r��5iv�` ܳ�=�8�#��2��A�G����J����	�}���EH�,_��6㨍�6�2s����W���Ҳ_˟\s��/�Đ��q�5b����h�y��[C=���uF�$�{��{���4t �x��A7n�"�����rڊ��b�mTXΤ��{Pއ�GK��+���w��e�w&�D�1�\�ή��	x��qRO�#
<�c5�o�z��I%P��i���Rc�%�8zտ%
N��� w�h?e��t��!z�nI���Aެ�����_O�gB� -UZoRT�?�����H����_��x��_�lH�_W�LZr�F�8ޏRi�Wr=�G��Gc{*^)��O=]+]�:���#2�/p���Ne~ؠkc����w/�ōVI �^|[�Z��z��8�#J����$"�a�h�C����yl�߇~fҌ��z{��{܏	�h�-_TDM�/��͹��M��?jh���+]/���u�>
[x��UH=%�$�U7q��@+5i.ru�迾��/�۝9���E}�w�3P�~cǲ���W�t�Տ�瓺\��u�4�\��jO���A.�6x���ٖx/���>�[�P���=塦`)���/�v:#�)?���y��k�95,�/�`Q�3�Uw��%O�����D�8�*��t8�3@�3#�ds�d���S��;�eZU�˼q�W�k�v�2��,R��Zo=9#Ra����`B��e���w�Oצ�7������:��f�)���d
��Sw��DH���y��F͋�-��t�W-s~�]�!�s�z1�yN����OLX�9IvPi+���#����:�>*���˨�D��)	�g��Rk`j�l��-)����joo�W�8_#ٿN���hr.�>_r\��u�͔�[:��5����.�<�!�r��dy"H�]��[V�C�Z�r~����e��[JGN�J��6	��)g�4�q���4�>4=��mmOӎ�Ϝ>x��#��z)7ӑ�LM>�w��]��A���:ڿh:M	Y�A	�u�%�C	sn��:���r���<���f��^:eQ���)4z/�@�9^�@=R��=�<��%���K4WF%Ϊ�P~��������˷���C��z/��˼�Jœx�jWV+&E
F��ZRKB%򑤾J�qǵEI,4躍WP$������`E```��й,��Ӛ+��C˯N?�o����6��+wY���g|<̊��	;S��&��9����n�0���{CX[B!�	'��X��U� ���'ÔMo��ɊZ31�цHN쓯I;t�/�!4r�6��º+c�"�����$-VJ�H���_j$p>[�g/|�Hҡhҡ|󳚉ڏ�E�e[��h*�jT�4�M#4�������'�brOO"F�(S����s�����]^|L�I-|��SH�����Ix�2E��2E{ �*N�[����2W]0�caR��媓޸�|��I���͹^�h�0���#�[S�tJ���$�6#N���?-�ǝ�����ؼ[�zi���c��2�&4[��ue�'�	�^��(���@��Ni�}����j���3�k7+�읰�D�P�r�Ι��T���Ċ8��!'��c�W�����I�פ��1���	 �����b���Y��a}إg{�mk����M]Q�g�A`E���������<C.��E):A]6��`�)��H|LޯnDc��ϋ�vg���OTdM�l��cJޅ	�_����q8��f}�3�H�+抴-�Oc�"��ər���o��,�?��J�D
���U���
}�{bf٪wW���Q���yo��\���U����"�����^h��|gdW�$|�~�/���Ʀ��a%�T���Ʉ��ir-~q�$�e�m�t
V�\����V�>kFP!2�{a�@�B�C�5�K����K��`Y��>�����S�w�wo�a%	�b��Ä&k2��2�����5���o�H�P ".S7�<��&�R���O�`#[���y��&*(�K��6	̹���.��L��d]�o��e�z�X�@�/�,�3HE�ʍP���$v\�CR]>~�)_��mBW�Kn���aA�E�qZ���w����L�G�3�{�C�A�o\+R�����q`&�'�%>6�Kؕr��IN�ZR<�J+���4�窀� ����9N&R�{��}]��06�d2�{�V�X��nA��T���zf��$�y��҆�UAO��G1 �c�S�$Ӟp]K�ߣ�����q5�!�<}��'� �&5�k�2�/�R�{��������N�D��R��'�c'cz4g�A�i���Ex�ű_lt��5�3p�g��T�u���mj�W��Ƅq��▽��o3�gR�q���
��m�N����{�ڽ�7�5�P24s���~�<�rw��E\_�1�Y\�W(���xM�Y�U1S5�"��N����Ǝ=�`�'S=�$����%C�>���*A޵X�@IaG
��ҽ.��H�3�.��M7��J���!��V�d��*$�j6�v��Pڕ<��S`�6� 4G�j�rK�E��%8A+xz�p���c`�:��� �/���x��UW���+w���4fżS�#gQ�ks��i����-��%�+�����?�2���+�	�q�H��W�'�cc^�+T�<s,��,�V�%�z?I�1X���a[��ABB1��"d�v�����^�c��IZ%cl���0,6	=��3�e�w��A*Q�O�
~�����S���� 0lͷZL͑;���lZ|���2�&�uh����dύ��A�����O�T�q�'KϺ�0M�AԯƠb��f+iҷcV�"6�f��IS����em����6��:�����^q�n�Q���`�y_��ڸ̖�h�� č���������O�5�"T���G�w���_a��0�Ҟ�k�D�j?��qt�(�O�A�-� &YsB�c�O�
,k�t�h�H9����آ��2�wc��ѥk�ИյhA��JcE�c�%�K����ح����;|�'^s��[�nЊs�խj0�X�%A>�u�$�=��NX2���cØ �g���l�tK� �^�cd_,�>f`�X'&���UR��^!Uݣ)g,�wlU�[k�zD��`���L�C`�d���vƊ}_��4��� ����=�M�ɪ�R�Br+��`�ɷ����U��4"{�ٻNr�V7�A�"��-JO:�������`���9pH ���W���_[����1V>�"��8����"�Av���;E���kAڋ��#7�:تJ$���Ӿ�O�ߌ�!Ѻ7E����N*s��r�yQm׽@�� F��\�,r:�����!�-���1֘�Ťr�SW��j�=rn��Z7����  �(R�ڣ ʲtn�������N�C!5Y�Y�'T�����0ְVs���ifk)3�"�538���/��-g��J+�^��`��Dz@�!�Ï�D�e�G�$��&sʏ7�	��@��j7���J���{��5��_~{��q���O�E���g6T��\Z"��65�����Ba�B��#c _D�n���yb�#aSi���ƿ,�6�Wv�V�)�m�Mg/gE-p]9����@������

+) �e����ΜleK4>�d4��V,����8��Zuc���)�6���T�?v\���h��:^\NH/�����q\��f̩\E�k���-߀r�$t+�i�ϸh���N�U	�"��K�`yQJ�[񬁰�bqA�1iw_ŵ����G��u`p[]�!�P��^��ZN��I�o�Zޓ��֓��ˉ_�n��Ġd/�)�n3ە�����E�8\����)�e���G��]3��m�P��>�*�H�瞧F���j���H��_����}_Hlx��'�ro@���ֺ�ag�[Q�-�C�X�J�Y��S�wȨǊL���v���h�f �!#d,O��ob!�?k�CM�Vu��Px@	d�h6r� ���K8�60f�����>q7�P��k�j�ݥ<�OL{�"i�Gq��Ñ=��Z�Y�῏H/����0E��B�l�	�]�m+'����������Ϥ��/��g7ω�5��*X'��2Nr� ���2�DǓV��;Z.-Ua/����<����J�
�Ŧ�j������ ]�=�(����k�M�vϩ �a�V��+(ۋ�K���U�A���� S��Fxa,�e���˔�	-1u�GRC(sl �m�TCQI���97�����10�rk�ɞ1����&!�Z�X�ɓ�RU6{�:U�F�ݽ	�rV%�!"<�K�W����@���j���H��	o}���tq����7��l�(9��H8e��98&��{&`�"�&}���/9E<tGBLC����r�l��.':�ǆ!O.�ߝ��� ��u�X�bDٴ,6R�Cm�^���n��/A��Xļ>x�yF�򺓾�� .��\lm��]�0�5D����n�t5��@
���)�s�*��v�bN'��[�����I��ծ��6QA69,jO�e:{��V���e����4��lP��F���6&�|ǡ{ "h�ćF�X&(�&��H���䲓qX2�!HI�읒⽖(k�[�ox�}i}Ӆ[�4��Ɓ���$.(���	�y��=S]�Tz��ҟh���n7#B��MsLdx�����{��E�u�uD̈bru��}�<�.��?��So�Jj�{����2��U�ᣊ��<����J�"~]�e�<ۙ�M`�̣�-���E���ڧ���z���)�� ��%Wm��ɰ��� ��E�j�π籠Wfm���.�"���gՊ��Wʒ�<y#��C5���hw��l�A�#���0�c���!$�V6#`����M
9���{��"�|W�*��zߓz	�}�`�X�'�̜e�dk�����I��Z�|y��+��WZ����ld�����bR��!@��~�n�c�3|�� ;=Yv��u�@������K�!A;�q��I��[��'�e�N��[|v4���}�5
W�/���|�7����F2�u>�T軕r*&<�SA��뻾�n�~9}�+�jq+�$�ˠm<�zZ�yҦ�s��s;=2��=�"���a��x�x�8f�b^��q����C��X�~��L�nC@���&�m�raZ*�]�Ö�o���_�œ��W�]��p�}�˫x�eM-�[��m����6�9_\�5�#In"?�\��ՙu\�R��c�k�(V-�v+�̰��Vaw��w�XL�G-���hK���-;;aB�bm�z�GR%qZx���ފ�ot����Qgm���=*�%�T��!6�vg�A0h�<2f��4�~n��;2��cPa[Lz;���a�����Z̙AW�<��|��iq���v���"���/U���+0˵�������yʦ�����e`J�u�O'Xd1{E͙bf�m���j�#�+������r�]OW�ٹ��I^w�d!Fv�j��GBV�C$��#9�8T4݊�$!�F��e���<���mP�-Щ�_g�&���.t{v����v�7�{j�i���6�~��]h ,5�5��+V6�$���)G���<�M�}�;ςk�9)�U�^xj��m�uE�q?ui��ލ�|���g��i5�]����ݮ85#ұT6��[do�g~��Ƨ�>�f0��nsU����v�/f0y�\CA���c`X�~ �T��#ŝ=lK'�.����;,�'���]�%[��{{�~s�#��� ��]/�aU����$QL�/��b_�<�"#/�Szf��gh%�ha�W�&�ϬO�C��#'��k��!�$�f5��-�E�����h��.�ZQ�b�6�v��ťqr�l��G���n���љ�]᭴U.�>�_c1�ٜ�e���@kAgy��|V�,�̖�B�E��z�>OVչ�r���~y&⟓�mh�%�r�`���
��]=_ �<4D�_Q��o�%�	�`�g�oR��^8�*@�n�������P�@`��`?�y�@}����":�|��p�MʾbN|U�n6�9�Щ��F�;��e��]�K�ΔE��_��\����==v[y����	S�h�1�*��ռ�kP�'\c�
`���D��L�g�~{� ��Չ�Ld�٤Td��s@��0���|���u�t�UZ
��;=�J��o���qd)��1�S[�T�ӳQ"��5+7`o�Qt9~V$՚b������{d�J?���}�+.->G�	HRh�6L�G$����W��raJ�ޠ3Ow��]���⾅N��b����Ƃ�j�X��7�i�vΖ�;����z���h8`�7�sqW�7��L�TT�	��57T�!���-]x|fߞ��c��ȦI�,�YA�&cC0���:H����=�wS�O��b�+zD�U|3- zI?�JR�����2xv<�~��^3�1��S/"�=za�����"g$ǭ�s�/��安j�2m|�w�i���/U�?���7�\��=��L�׸Yy�Ze-z��̪��������,4Ϙ�=�]��fL@g?��S��c8��Զ*�4|K��5�}/7D|%ʲ����"���ژ`U�[�[|hC-��vv��~����d;�+S���\_��@���	��-�6�D<y�r��,�o�:���v���۠���1�g���!���:�M�9���zl�A�]�L�.4�ѸK8>��GK��*F�n��	��z��D�:��k���_!V�ø�G�i��0����Bf_0�L�m���� ���P�VfB��ǈ���E&]�OO�����e��zsH�Zy�g؏�Ŕ6����g��0@Oè�M@��iJ�t��4	'�F~�1ԑgo�ko�
����Mn���h����@��� h\�� ���V����t��iqE�!����#��*q?M%��Ƌ�h/����J;���Hk�&o�xz2�3򁺆1h�3tsz�#��nl���xWO�/r�Ϧu&	m�q�?q{�Gu�������!�]6�A��b�0x??��'����SPZ�$�"�xN���0�e
c��d���� �|7��wKɻb�i�>�;����Z��	���L��#�5W��8��_��]h�J�֜xX��z%�Ɋ���c��� d��7�����BQ��z��ٓv,�sPI��ٲ�ݱ���mz�ic������
�]1`�=�k�/U���7G����xAkA<w������{~���5��� /N,�f�����EH��-�l�3��m����ޡ��a��X����Mt���ɱS�˱�*�l���;���0���F���YUb�pk�~�r�8��_��EսV�����K�m���&��`bG&&f�ݡs}�:־q�0?�1�-�^\z�-�@�?6��?���E�\*��#;��e{Ϛ��{�3HCs{�k��Q�j��>f�P@6�&ps��j��v(atc{A�lZ��l�5��`��H�����v\uA�h�5�'���]�؋��\��h��Xe���D��,f��r��K1��ZY��4L¿Ѽ+	{%���O��n�Ӯ
ԁ�*W7n��C7b�Li����+�-8a��m��ŏX2�[�Q��6,p�� fEEɥ���A�s��
e	!;��m�ڱ�Z>R	N�L�#��	!ʮ})�Aۍl%���'�\��a��t�.;$��!�La�����po�YF���߻hƵtA��m
y�V�b��4����Cto�@��T"C}��Ѕe�R\}��J���8p����AL&����e�4��q���1n-�}ƀ��L:1	J�
k��^�/9k'���I ����" IR-9!�]ר��a�{����N�� �b��Ԇ��63��{����)�i��Id�(���x3[D��l�h7�
K�rdw�\`�q��Vl|��U6HڟV0U�����O�Iq3+֔=�l����8��LsX$nR<����� 2�G�W�6w�c(����	�q)���ݩe�%DaE�!{����Ȟ	REX���H*��EbI��3�#�'�08�,��z��o�Z�w����^���s{�s�ȷ��ұL�4�7�u�8��
������R,�sP���8��x��6�����>�L�D�~�΁�0��d���,�b'�����@���jP���'%?F۹p`)���	�(A�=�#�vמ���9��6�����{�8d�_�,*>5��x�jM�-�����;����C��F�0�!�:�z�Vv�_������%�]/4�X+��gSu�YDW~9��}0T��4���pQ��<��.V{S�&��1���a����&!�&3�qxX�̟�q���-"��1"�����Q��#����wzx�g�q�����O_���&X*��M�0�T�,�lի�_��=C-�
?�����1�[٘�j���*��Lߋ8���g����e�9.�6]�� �_�pX����J�Ƨ����d�g�'p]�'��w���E�ܯ��R�����y�D?Mo���X��>�Il�P�O�����}�/�oK�bIV��i�_۠}�?t	Th�i�5�|m��P+�P煩%{-�����haM��ݸA9�"C6h/}G�$=" ɪ��=�Uy"�>����!�a(1�HJ�Ɵ6Ъ��lDa�]��w�P�tx�`G��x�f�y�X��#êT
�������+�����&�B�SO���f���8��#~m�T|f+X�TdK���o�Ƿu+��Q#��"�������[[f#��֪l��X���@ N)c�Lr4"��ƄaLo��� 2�E%����(�e���q�'�s-p��7�ci��,��n��sd�q�g�풭�����7�����VЀr/w>�O�6�tn|w�P�#e�]kN��')� iZR�ZG�9�g�~�`̻� 9������juI�+Rrʃ3ҼecEij
cŀ���H�1��J�*g���uͰu%��x]U�6��-r�a���6��zex���ï�жdXq��v�q�v��:q�Ͽ�~jC�|�X��Q��|��,U� ��>����2�Wz�O����.�\�F��QA[��!�vR�J��v������j���Y̊�Ӄ��в���u�`��9?]("�GN*��P\���rrIᰅ��Y;�˂�k��m�G�Z�L�x��Z�� ���=�陡%v��un��>��Mk;��E�q[�"� �2ѵ�˂�Dں��Q�VP�q��.��E�&�ȠSML�	y��n��s���"U�&f�8
���}�:�^\c
��\�+9UL7����cn�^^7���}K�k(��*���zl]6��8�]y�7��~ݥ/p���A��@W���y��:�0ΟC���T��=�dk�**�Q�~�L1����n(��ƃqK��tެ�Y��T��e�0�JU��Jy����H�ɷkL4Hk��o�1����к���Xm���-�8�0��	L�?S���2��8�ק"Q�B���#�$��n]��)$R;��{}l�8N�FbR�!렓D�\��%ȆK��`#a��6oy!��"M�.�h_�f��� ��\r�&�t���;�`K8u����x$q/��<�}J����L�1lJ�����ԱP]�Ť�5�Ϊ�h��Yn�Eo�=\�Í�F��1�*凿e�ч6��ƜY�v��W�U�Ϭ�z�i/ٰ6%��f�9un��>�s�nm�����p&�%�tڶ�Zg��b|�N�|���.p��������HJ.J�����ob9�����
�jb�#K�rKҿ��ab�m�>�=��e˩��,j"/ ���3G�dUx����0����ۼ�9�7�><�v�_v����*י-� W�����X=�/+������fh��O��3�tr��ޏ���j��E����A�S{W����a��ن�^�9��om���^4�Pj%@Ӳ3a�U���ߋ�ƨ@�Ywr�><Ue�qwvɮF����E�ѳ����S>�쨾p���p/3��v[���ib={�˜�W���?�c2�8Ы�˗��qo?��:������I����v�
� _�s�`X��3����Q���"iG:���0b�w�`&F�ρ^������w,�V7큸��%|�"�Ƶ ޒ�"D���X���`:��V�4�ﱫ�=8:�9�pW0I��8(w��:�vNh�caRk+%�b����H��~��/}��,hb�e
�)�Ng��H=���7�;���`��"!�U
��G�~L=��O3�Ԭ+>b^o"��o�%�ù�1�@U�O��(M��H�U�cW8���Gɂw	 ��q����S�����]��/~e��
��Hc����-����!i���'���-�v~��+�˔+zlGi��xU�r��ػ�K�$$��l~}aK�0p��N�R-�����Z�A/D�1����6�K\�<�ţ�'��w�Jg��K�Ev��:X"��9�9�z�.R���Z�V���o�눹�������nh'��2r~���]����Cb��q|do��1���$˖�\y�dHצ���ػ(d�u�t*��~zcCt��d�С�LP?��̙G�e1�(�A�}��ga�h�oðk
�x.nQ+���L�����C���&��0�
�N����V��������S;��r�	c�u�쩡�P���"Q����lm24g��gsv_��,���?�Ô��<�o%�����ť��6���{xr�ѵD�X�����%F#�Zepx�#2���$�NZ�IX�e5�lIn.8���=b*���M*o/���0]�lY)�rG�d���*�4�-�G��o��\�4l�ګ�y���T���.��+<�A���K?��r��'� к��/ �W�^~�@����^��Ew�ZG0J�;����"Uh=���4��;�!?0�8ҴO��4M����i��7фG���ڲ�˭����Z�D�m�b��څ'0�*��ÍrЇpк�hR���_vg@�4�WA�x-Ƴ�Ѕ�~*evf��?��k�0�(�<͒�8�"*��~�S x �zil����,�=���!x�:��;��,r`�s�AD6g��@���{gT�}�ʪ�;�w4��4����|=��]�ƵW�����i�͇ͨR��7�?$�%�v��$�5'!��q,�m�d-w��ͨ`�&��QS�g�y������½⇦�w����	V[Ϧ,؋͌l�|����_\��sl��L6P���S��s�&�T&&����T����l7�>K;�+�#O1����-(	����Q�*���p?���؁��>��^�ֈ�ȳJ�|�ĄkV�)���\0aD�$�o�~!C4�zSf�9j�_���Oi�
�+���)��ڤ�P<$��}����9�������F��c#��L��m݇����A+�ݡ�iUeo!�u*P
��@Z���fl�"B���1 ����[ã�����PMU��m}0��:����kԮ2�م�֩�nf���@�F؃���8~��U��K�R�7ՙGoe(4�e���i�@��F�}�<�<�k�"'�@��;�ڰ:�!.\�ŝ�����Q�:$��x[Ur��&U9�$�Z�Y��A�����a)�#�]U�6\Dz}4&���a"1��Nu�&�`���Ŗ��w8���l��6w�^W�i�4V�h`G/V�&�_�L|�_R�M�[�[~dY��^n)�9 
$V��2-o;�T=U�P\h���c$Ԏ&��>	��PLo�fy�����9dl��Bٙ�z���4C1u��e� {{���jNITL�t��IP�o��F�� S���5h�^��0U.�G��&-��A�~TM�Z�f'W�P��*d��_�mH~�1��w�e�l_O���S0_FI'{u^D���0���H�k��ي7r����
��>N<}H�Q$�<�n�[|p�__�H���y �MҞ�r���z��A�ˮu|���k>�̥��fZ�`@��N̼����~V��7�W����ʿ����	�O2ãގ���f�T�@������j�;��y�Q��4X&�MZ��#����Ӊ:��:��Z�o-������ s�pYw���&5��I�RM��������|�����H0�V(n��n��:Z�E�lRǆ^�7 /`�e|�*0��0�eI����qڽN���uÞ�#W�	���G�
/i��h�2���vè���о��Ծl�7a5A���D�P�
ZP��W �}-i��hA�̪�042��e��k+�ɬ}Q��|\p�4.\�aֿ'����$4��&9�GAsL�A�ʹ�QK��BZ�B������ȴ.�z^��1��;^��	k����⫼��i��J�m�`�ڛ�~�bM/]c)��ջӒ� �	��;�X��L��=.�Lt���pK��;�I�L��l���bu��{��LcK�A-��|Sx0�^NJ�×1����\!R�j-�P�X�)M�P��:X�o�1tOXh>)3,� $��45X<�m���h�k�Qvy��ԛ��\�~�^m��3X��6�t]���Vn�����YUT��1/�?�n���2�~eׂ�Lj����=�}-��ʯ6�~��[��3� ۔�����R��������e��V\u�� 2��͕�߼Z$%m�L�KR�c�Q�(��y���Qv�'eG;>bc�>�ˇu�s�4+�����������{�)+�P����Ϸ�W����έ�z���>A�6��պaGd��@���oj�^���0<	M����(�����3��I����k毜1-�z����G��~S/�/��տo�N8���χ�x�ƪۈ�|��r8�	=ܚ��	���4��c&��p[�ZX���k�ў���e^F���	����v�6��6:��[yFl���:�A��F
N~EC�I��uz�ݛ�<���a�-��.^<o��/�u�{Ӥ�u���So��Ŕ��F޸�AR�z	1������S5��IīV������k ��4���!�����AEe>��[���p#h�/w�q�����2��M���ot��;ǌיpD�>���\d�ϙ�&�o�LS*K�WX� �t1�-�3u&�w�Z�5�Pt���.?u-+-����W�E�	zT�Ei�R3FD9;	���/_eHx�+5F�-��!��,r��p��<�p����3h2��E�>���34i��a�ݥcTY�o���������������=n.��/["�E�I��jR5�kÚ+�{��^�p�CŖW\d�v�[�k�,��BmRR��-�qҸ�����c�cUچ��ͱ�
{�L���:��
c�'����\��	ʸ��������^���o�G% ���O�5E9E��z�	�������^ ����d��~�1�m͑�X�[�p
SXb�]�4�
��
��&����d�y�(����
q�����aU.I�S/i�5��G6��**�G2>�M/񝆆Tf���Gd���X���#��yxz2Z���h�� ��g�Ȥ�_0��LiH�`��yV��[5k�A�;[��e�G@�e�2A��F��_�M\c�B����y�TEF�a�ڏ�UB~n�����c�����2Ŷ
vd�R�H"i�]�`�`��ۓA$�rs����o�P����x���L�|��^��4Q��d��f�!���aVY��	oዖ�n�}����~A��-�28*e�U{͑��TZ��sKnB���r=���Fw����7������.��!1�k����a6]������,�R��9+B�p�;�ޫ̵?���e��K�Q+w�]j��W�ff���i��3j׭R�+������%֮���?�W���}��.��T�Pa�&u��8�4J ��u����sF��u�p⛃T�t9�Bb�Kc)�7IY�bpﻧ�Gsh"��٫S���S����.꟟�k��kAI��G�]� YK��U�a���lO%L�����^ȷӤ`��� eo��֩�M�D��H<?���J������dA��6�nM�XYe��@,s���J���+����ߘ�E ���Q�sRM䖜c��Ŀs�y�J@�l�'#�fR�|�h����S�����Δ�k�7aI�����EA��b�ΰ��y��=U����;p�^Sdh�RQ~!��CK��K��_xv���)x.��)p�%<�}c��"���Z9�+y�E�R�1&S�<{������o�����)��[��tkSŽ	l쀛$��w(w~}�C�����ר1��Ѣ�ߘ���)&׵L'Ғ<�7YU���i-�� c��'DPT�E�u�s���X!���VO���^|��,Ja��g�D�ׇW�XV��O�Y%M�!}A\���6�����QF��[�=�ա��q"�o�D�hn�?�[�Y��/��`�w����&�0��- ��M�'�L��Ė����:�^�4d����ʼr��b�Ԅ`C���Yu� ��K��ޖ��M@��ܾ����}]u�7�LvU�IjJ�J��<E���3����"�j�{� �����/A�o&}�Y C����-t��E�C�|���W$δ���]�EA��\�׺�ݯ�3.�cv5�����_=�|"�1.�B�N�(����C0WT~{���U��������=�T璈��+i�~ի��p^<���`�Fx=���?Nr5_?k�����<&F��m��f&&�Dk;���Hj{���?;����F�o�q��Չ^j~�H�7���"�Ͼ8dNs|/����<{��(���,��K���י�&�O�����g�=̦ا�ޒ+�Z��_��PO�9/���\]�����\�KgY ]3E#1x.V+E��hՏ!��yX�����5�?b'�L�+����o6�Ki@F�B�BB�W3y��Gj����Q���w�~��[}^#]�v�q�o.�����oxY���!w���m�4k�1�\���N�s�ȸ���Y&�y��Y&?�����NBߏ�k�|��8��R��ȧ4n�:�i�zm�Q}�LBR{� EE2�@?5p��������ne�t�t	�H�tJ�twIwݭHww�C#�t���� �}��ܳ���_��z{��y~��"���J.��9t��ܪ<M�1h���_��7�W��)}N^�'�^"��S����XCV��@
�hf�mKt���w��%�
t�w<���k����Dኊ�P@�\E�h����w�C}����n�ܟȌ�	��عg�$'&�&!�
� ��]�C�Ê�k+�VzI����{Y���c;0V1pQ�Y�*��˺�}�O^��e��!~VHL^�p��X�������� =nnF�"�\*H�l�/��̔�NEu���坔r��[�[âu��/MY�_����qTu����s����+r6�mG9���p��/a<�ņ�ey�G��\�2Ͷ砹�F�dfeJE��t��y�G	xbXvM�Aš��+η9&��/���~Ѹ/�����؍� z��g]�6G�< |��&���CQ��{_83�z΂4#rj�WR������և�N��ֳS�V<Q��[�5�*��F�f�U4��R� ��/ۃ����]�p �J+G��� �ڭtg���敬�w�T�]��T�yXU��5iM���Z�v�qg���vvs���Z���6n��4���}�>d��xx|�m�P~:\�TWK6��>iu���1�G�V2��c>���rj����S�����$�K>�%����
��0�Ŭ�0��qV������j�Rh�����M5�;vp��R��d(���a�b��1�5(����9n��Q�\x���X�?�l��$|r��
�S���H��}��n��j@}_Ǖ@����j��shLE�bl��|P΃S�ùW���(:H���*̰����rc	���X�d1S��9�vrr��gg��mtr˻�1�e�����Z&�"��f㾉IXA�F����p�ס�h�=L�D�Ґq%7v*���`�f7�b��=A��A�)	����ȇ}����u��������z��8�-�}����z�c�]�t�s���ͯ=��gP��r-�\�y�g���>�l�W���#W�v#Dߊdd.�;o��Fd��>��X�R��] ��|w������RPogi�����nz�lͽW'�`'O!(�+oφ|Y�`�N������p��2����T8u�Kǒ�qg�v�j�fT�@5�.��hkC~Q8g>	�t��w+���4V+���"(��p�����K�����Z���ϗ�p�����_���юe����`��eI �]�ar'Y���Fi��͈��i'bE���X��L7����Uۍc.�!�A�ĵd�g�q��-�"�*�|{qu��$���m/�t�c�s���=U#;��J@��Yp_��[�0q�1R���C R	�%y���9�kB�j�!��g�ǫ�	�١�bU
ǹe\���J�7UUy�tS�C�w=ϤwK���&�O��qC�U��R��\/��!e5�nB�9��YA����:���u����(bi}¤�U�hf�//��\]�cT�/�9Y�uh�,D�%!ͧ��h��_�tX��^���O!�A@��kղE��!�Ѥ>��#������z��T((��_�J�;_m�V�j�;{LZ<��`�t4���jXgv�C �b4U+UD�k��X�z��̷��<�.�&�K������CS�u��e��a�	�[q'��c��R&��1в��jEz�K�IK�ÿS�1F����}�)��;ͽ��c�mWx� �R�i�K�K|l�����^4?G�����F�F3�&��E�|���hd��J�w���I7M#���vxj,�m=, VTV�*:$�i�(��b���Mg��(@6X%�
���:����~�xz�ǹ�&2�� �_7�wx�����5��#�Cu8���o�;���g!��
;ɑ��ջ'	�J3����"�_�@9\���\���z|��<��W���u���k��U�����؁�t@���_\�N�~>m�3j���M�'��H��{���iyݻ��J@ %����p����=����'W�2w�I�V�)'�ws�'N�	��6�d�!�ќ�g�a����r��Ϋ��9�}�ޫ�&�w+Z;g�>��3j����K��;���J'j�OO����(-vP(~�^���g�@��/��t��0g3]�
����?ҳG��oo8�	G0��|��S���rMQ��s�6?��o⹆�&���p��@&X%����s��Xj�ߚk���G�r�Rb��x��e\d.<���xy��ý��"���t�^���Ûo�O�N��=��paK/ӽ؄~LV8�g1��U߷4�R�̈3�X{H.��o}�VjV6���Q�rP��O>�	�Z�>���/�b�x��ƞ�]4�W���/k�B�R�i�i��s��(v�_���܊��*�S�������seʰ]ֳ#�_?�CJDr�b�"h�8�Z����`GU\��֎P�G��=K�%j�L�@����?	>M������Nb�4]Ƴ��*R1�9.��؞��YM����_95�S�y5�b����~0�+T��ޞ7���nn6���1oO�5Ln6m!�C���N����j����'���&�=�����4��Lh�"n���U�5�<��A�<�g<Q��Q�e�V��~v7��o��ZTv�y���k�"}��^垆�ֳ�I�vaŴhl l����g�2ڋ5_vɁ��*��&�����Rf�؞i�.��\���p�i��!����㣋����U_+X�ޣ�X4�ިDB��'�Zh�z�����C�\����)��E��>v�wW�֏�u$t�M�<�F�'���!����(�l:�����cE_�׾SF���jK�X��Be��B���n���MB�ju�)j|?\U���i��묧�"]��)
��I�t�����u� x��k�/E6�@���C��ܨa'�{���N���z�� +����L��1�y��z�� ���>Q��Fk�ϧ+x}�쓹���A|C�:z����М�]pf�Y}�{��x���'��Ķ��c�2!�����w����8���
:�+m��\Hb<���M���4��{tb�����z�7��8�t.�xiɥ=TZ�2� ?�s�+��:2�8�s>��$�0GM�M��_ZSQ�k�e�"�ewX�G�r�r���!w�.�s-��.��j�^{/��ܸ��ʺ�֦�A$�V���r��4ܚ�BA��"��{E�U.4ȓ�F?/����S���A:���_�5ْ���<�-�jh.?'x)h��o��DV>9Zl+����^������1�� )4Z��3��l�/��*kz}�ʫ�=H�$���2��k�Y���%�N��;5�S�}�>�h/ �'��W=��űt-9 i+�ᇖ<�����W�q����NF�P/ �A�Do�=(�V�SK�SD�Gr��]�������������,=��Bk���Cz-j|�[)9�ۅ�}��:	G�CW��!��ˆ��*z�U��b�³<��َ�#�������Gq����Cip%_[�(R�]~	����V�
��*������#�R��p޷���Z������RO��{���0����.D�k]me�E�Fy�V_�e�"ŧz�����8�D@[��k�&lQ�����B�Z�����j'�aϿ�z�7y�MZ��5��*5�V���-<}�#����F>%}'�=ŏo98��8�	59�v�O�x�j�Dz�S��A�]Y�	{�T�7d�����g7��U�,���>���
�"�b�P�J�lLq"߆�i�UO�����M��h6����H�!���O*��U��ҲC{E�����������O�PU*�Ul�}�}G^jH��6��*���Hz�	��m�m{ 
\b_��k�u��_�:��b��=UTص>e �	<�\
w�vL��1�-0�h+>nK�l۸�^����ݱ;�|`@}0�C�!pnIk��9�st:�c��D�������D��1�K��QoK=�e�'���Ui��]$��Z�rI�)��z77���� U�!�{S�}d�l=�����`�E��.�����x��\q��I��B��9��w4nم��"K�v�淋f4\Ѫb��	A�q�_4��H���bO�l�Tᇗ�b�w\a::ܤ2�8mױ�^������+`+5��n��_[���jA�qh��
�I��E9�M0cJ`2��r��Ph� �V���Q3s�,w5������V/o�D�?yh����Ӿ_����-N�� ��U��r{8�Ŋ�A���Rg�ջ�>zA��(pew=x��.�"�{?cd&ǯa*ΰ�cnF���WTdd:�&��>��+*v�S�,���|����V�w�I�u�W ��\\�3ױP�$W�ݮhǧ#N�hl��7����^�A�����Q��eN4�Dϯ����Q�1��7���g�=����pyYb|9��d�@�5*n��<2���{JmIra�7�����u�hV��:٫����8$�B��O��+����N|/�˛w�I�%���e[�.�8��wj}�p.c�K�#�Z�Gl똞���O�ܵW�~p,�y���2%�e��a_�%}L��^�N��6�����"��S�t��Ϛ��JPd�|%9R�����ܼM�_p����Z( �@t��5S���k#Amh�Z�éB��ONI�`������K��a�<�H7��z�kQ��"���6"D$v"�h���8��K]���	�Y�w��&JV�=R�*�F7�@�lR����4�3O���R�]�ɋ��-��}]"���l�A�+���~9�O@�7�'�8�!��ٞ�V9���q2�+��u�m��n|��c�O�0J�w$鳑V�v������$>��|��H%�ܓa0����G6�2�.��͵��/�6���8�R`0vK��z/}t����X���ͣP?� ���䜀�m�n��ws-��|�� �h�݄bΝ���5�xw���o�Ll�6�L�4F�:@A}>�q<����לd̒�ٮ������s�g�cfF�Z��5�$Z���`� z�����vHr���!ad �w4�*��0��q�e#Z�z�r���y��|H��N���Q��=()�/�l�Ժ�n.����5x��p�H���i5}�C4S������qRR�M������VO!:��/丳�s�G����Q�g��\���k9f1�*�Z\��p�����w�<
���Y�R�f�n����C��_8��}ER�.<ݨˤ��F��{ٹZG�<�D^��P����@�8����:T��v��] ��Y���Y1Geg���X����X�����������p�1���E�
�}޼���wHA��p��C6�z~����槦)��2��>0�*�xy9�������g��'��C �)q�h/�sM1gc��b��q�֔H뇊z��,�~9���8R���w�6�<� /"wx{��g}�1��FY~�ta�ڶ��(�d&�dFm�_=�-�،Il�3뼻��J]_}�h�Tvp������K��kYXȽ�8'pl���Yu��w�Mfq�
pE�m^�/������3ǧǷԾ�t�-ѹh����S\NT�;R�U��&�����#%_�\��?�\�5*��{��aK(���G�ݳ9YVy��]�n4�Y�[82�跨��Z0��y�����i��p���t9�C47���p,4�����t��I�f#T:�e���]���6��Mjw�G�1f�Q!�Y���[:��J�̴�؝،���5IBZ�Ke�:X����PK�W��<��я�(d=&����|�	���A����������^���X���#��3�D~~�����>�Of^��9�|tHe{�Ff]���N[fLT(Z�}���S��C��X<�Qbr�8Z&6� �LT1�/nz�6�b���^��3�WR������4n_����Q��k��Z�1R����R-�7_R4��a�k1�[�t���ܼQ-�콈�ɺ�q����H���4��?
�F��s,6��r)EJǍ�c��%���J}�$e��bC~y1:̘��@#++�kYZ�Ǭ��tWgmҤiP���M5��1AO��-���6�ܧBt�0�\��N���U*>#m�#��4�B�����������Oͯ�R}�a�7[�D�晳���H^��M\��R��E0x;[�\ǣ��_v^�ʡ�[B�Vc��Qk����x)�B�m���5���)6���
 Ճ�]VcO�v��>��)��`[c�M}���h�D'��c��\�S�;���yQ��J�L\����]9{�b���.������ LQ���J`#����T�2�S�ͪی4�2&����I���H
<bI����������g%K��6Cʻܹ�a.��|K����"��7mf���7_�]��b�|�@E�F��XN�}���Ndca�l��|�I�r2�Tq����[$��؂��������:�QD�(��aS��UJ�d0����x�)#���6�DgGGd�*��bc���\���\j����N�+�2��ͣo(u���QI�;B|Rw&O�;D)yif�q��Xv�����|�U��~lp�"�(Q{"��ι�W�9d���ޓaX���h�O4xZ%��'�[Ǡ_��Z�_�Q1�c��w&g�/}�q�m`��q:d�ET���3s
+�_S��`�����D��l�$�˦ꐀ��%�%�e;�0aK_G'�IU�@\���"*QV޾��j�^Z�y硫*H�����c��:HhWEy��;�V��a��}SS���L����!�{M���5ؗ쟶6��{\�>@��A���{��_\f��]X��)�6�tU.֎>��<�Z6�2����D���ۼxR�O �������G�C(�o����
���.�T�T���cJL��E����������2?O�M�W�v�6��6����I�(����fW��ST�DV����vDs(�B���m��H�;?�~���0�?�t/�XEK�B�cn��?5��u�Fb@h��z%��a^n��� �NbM���w.u�\a4^����'<NNtg�UX�~
���� ��i�vh���D��E(�Fo�X-���}����m�c��b����4�]�D��W���2�~ t	��)aP�~M�$&�cܻ!��X�9���@q~|o��v:7��XI��QQ��$�u��B�C��{�]%|(D�q	�	M�D���gdt����b��{b�(k��K#b�f%�fL%x��8�=Փ�� ؽ��׮P��;��q�Y�Y������
�1�M�+�3+�I�gɲ�ʚ�����pō��P��?q��_Ứ��S����Y����<�8�_�0��Ud��I��<q�;R���d[�ލ��$�L�co���QbS�׀n��~T�8 �j��f~�3x��媈����B�Yd��m��Ѐ�;���j��K���v���дГ�(v� � :c�7��Ja���x4��c���s���r��hr��\�n '$%�y"��,��Ş�
�j+|�X]Z�kA�Z2w`��횞�φd:�1��w�7փ	�W0DZ%�B��\Y�\uo�p
p�b�.��#F46Ʀ_^1����5�T�����L��y�j�k���;6��h��� �#!����654���}�O:�F.S��on��G]����J�{e��cY��M$H�%~H����8���k�ÿ����̇�OsE^���\'�o�Y��/{���z#l�AH�FK.�F�@����;�@<�����a"�nĞ�z��ݣ���*<�>�F��=1���#�xVG��p�����@�`kg�Z|:�x�*���ݚ�u�#�2��hJ���GRÃ>����-k�����J��ȕ8�5굎�Bq�/����i������l�N�ۙ+(��:��^8�fi����c����]/�D<�=�%�A�3��xx{ܸ�KïE��B_�Wȑ���Kѷ�'w�_"��'>����ԧ-���q���T�{�����6o�$N�x���S��3��[���?z?��V{"����<a��u
�%��P;��-����ͩ�"�b��R?��w:�.S0�xD��.|��y�5���9$��~d��0�Dt��7�`���=�DW�j���r_D��-+�o���W ��H'tg�6��*���q����x%�!bܗz0Ƌ-+(��S�}��^�����O������	�H�?񆄦�$A~8�=�g��Vr�-K5�g�v�a����.d�����Gl/��!����ha}N?ڧ�b�vO�{���6yG�0�ׯoauS8��t���v�$���b6�Z<,�Tׅ�Ћ�'v@�L�^|���3��c�fFͪ4�_�����$�i5�*�c����ܘ�Оr��&��'p�p]45��EG�E�oB���GS��������%g6�1Me��,uC���A��[[�V��n��P��R�Б>��6��^lx���x�4wd���bSE{��� Z����)�I�`��풒
�i��A��撡t��BzM[��k�8�O3B�
[1����-]r�#W^��7<�u&��	�s|/߃��$���
��#����Q�OS�X�'<��	���~.��ne�CW@�&��p��9Z?=MM$�W��eo�$r��Z��x�)��v�wB��J���DVfk ��M(QM����4��7�𰳚~D��Y�,�Q�C�N���-���}���1�'����z��v��6��7Oo�Y��nԙU��48^'t�w5F.i����eq�b`v�s[�����>z�Y囅1��y��/�$���L�r��߇��W01�4�c����=����{ O�u���s�lT��|��-w�)w�R����W����=�ί��]q{u�|�C.��mf�ꪪ�/�|��(Xo/�w���.�(���{@�tu���`,5��r(x>�6os+7PWl���c��As����rM�M���ht�D������%0����I��h<�m�r��[��D����� @��Ha�-����\�VO����&o���ܸ�m�����֞k�5�Ã%߅��v��s�DH �
���W��R��y�Qn�D��g^:�uL����ԁ	�N. ��9�`Ү
/!@�zU��-�z��ORx:�u��ˬᔬp�73b
8��F�V�i��w@�%]W�t�ĭ���j���ÖO
6�L������������4���G�SU��\�|Y����%%&��ݮ<����lݯ\��r%XK����7�B���5��d�� J�����ᣌA���O{�=��#BMuhu$�u������Y�oǃ�N�1�MpFY��&��!�?��r'Z<���66��6������b�6��n#=&;�Vh}�c��7���#�������^��MUl��e�m|�@��3p��zT	�Ok�J�`�j�Â��{	�c��R��Q	��Z�Շ����^���b[��3���Z�3���U�(qD�i����/��n�s|��f����`���7���-ϋQ��;>����O�2_t/?|�#�A�U<]H�r��x~FF�`����	@m�C��+;���4��<�,w�����K�4C� JL�c�ɰ�'��h���d�P�FA!���X�'�rs�H����V�,)����DA%��Ǟ��?��-�f-�8~���"r����k�4x������r͸ ��u�2zhO�C3{���<eJ�Q����������h]�M�|[[q�i�nm���#�G�l�SjǍ�/�'t:)R���ZU�y�ڠ X�M"����W_ ��<c�.ta"��� �6�����t>��?we#���o>-̠��$�`����t���p�z�1�qc����
QLA]}d��)y~\�vQ�,Tڍ{�1`��5�FoŤQW����ɗ�(�����,�++0cGC ��q�?[�:��@�p��V��	)"8�G��vC�u�n�7a/^D�Lq��{PdՑFfA�bw�X�#��)1e&�)���k�^[BZ��9&y��7�fK���zS�z6SEU���P�8y��t��C�����Ot��nE�{KJ����g/�%\0BԆ�n�%^G]/L�oR8�6�Ղ�c���8'�^V�m�3]_����xȮˮ-_%C4��G�?9-��.ex:f�$�E�����I�ӽ��'�"Cjh��b���l	u���ơʖ�ߖM�;O�W��u��!��R���m$"�愒�����N�*�.�����
81�6����s���1�gΨ/�Z?�5Ppft�y8�.7�uf�L@�?��آ0��e��щ��i_���,;{�J��&���m���mo\ß��E>�k�3����	���ʄ�oR�pu1h%9nv3�2x���bU��Ȳ*�O���H�������Q� F�3]2���{�G7%�G�n�}_����!}���7[ҭ
_���<��ͫ2kƱ��' �$<�Ez�7O�D?�g��eO0��:���@������������~o�J��I.��Fi��)1���'�2:!O���BHI�I��y�7�q��A��P���� f�{�m���~�^��@V;��T�P;����i�v�u:��:o$�@�ة�Os��S`%+c�w}7e3����zg�.��i�/�&Ae3.I���#ɹ��C���t��	�4A� ����_C;)}�sA��[��Mo=-[�Q�~��>͟fn��������Ө>��g;�t��n�H��+���תw�2�W9)�&����/�$�,T������Tܹ*�;g\ٜ�:]հ�|u0K�ġ�H�2��8�w�ة)4&u�����vgC����M;C'Q͌%�B{a��q�5&�nD�Ж��/�i��+�ؔ��=ժ����˩Ww�4�w0J��2�Vޕ�>���_2��6=U|b��~௱?��Y�9�_۰�q�q�C��\`�h��D���ZJs~���Ps(j&�kV��b��|���H��>��0��R|�^��?{.L�,�^"W�D�eW*~��DP�^�#��GX�Hc
��5b����&����R)���C��,woԑ����v�n����M��X3���:26���U��<�������L�������X�G��E,����k<��!����@�!�����Ī솵j�f�f���s�T#}T�㰅��rHu��D���3���~_h~�����K�r_,���С���$�X��P#����3^_��i����UO�|	�%/��vt��E�U����.�y�C�B�q���%ʥ.|��g7@�
/ޙC��p����WP�?�P�h��������Vr��	񪣝V I
���T��e�M��`tBL��kl�3��r9Ӷ�Q���&���@\w*����*H�+�i�����#�$��˂���W�(��:UT4ȼX�ݨ�V*M;��B�hF|��0S�*U��ഘs�_)�*�� ��v��]6��^}�+�����SK�n�Ɣ�dE�nc�e\++"��C'@A�� m:R���[**Jm�.8+�i'��B��X����Xk��_u�AO����8m9���W�Z�5��K���V<L���q��n�m����v��'�G�.�"W��2�"|h�Wj�F�:	�QS:)�@�t�����2B����o�j�A����7Ƨ'�f�,��j�at�B@�ƨ�.D"�H[N�<"��b�����_6�o�����HF�u�m��P�4G�fBo���NJ\�hH�Ѕ����RZ�G��/֦�����5���o:P)$}"����wzE�rQ���!�1�$�?�/v痁R2�+�A^��[?�X��[�R���܁s��R$��e�@�T�kl�5RH_�H8�/[�����âV�M �E|� v޶����5�7��Y���e�؆܀��*��QA���͆�i���W�4d`m%)	|���p��J5:�y�Ý[��-��d+pss�S�"��s���_U#2i�}�!���Z�w)�ncM�[�})p��>�-4kB��	79�Fj�R�1��>uu��iO"�-|&{Z��ɼ�q�n�[��R����8Q Vl�J����W��^�B)������vLת�Y��P'�Y��!�4��agu2%���[�SGg\d\t"�Ҫ|@��l�tR|Q�Yx"crk�㏅s��A��Adm\.щ��M�L�Y��d��Xq��7��G���rC�04KB�r7�J�5�� ��Ù���T��%��ͳ�����m
��c�
�`�k煳G�����
���9U�kVvW�z��e�1�*�q���[SWS�� b�8u��(˾�-�gx��H�\껯s�z�.��%��%�y<xѥn3������*c���htd��~��Dp��=� ���Ϳ�P�h��j��"��Y|{���������X������ߵ5$݁ӥ�A�vQO�X�ѫ�M��Vht63�U�L^z��(��#9�s�p;?}v:�P4����9��ue)���t.�6�{~a�.H�X�DW${�	����]C�����~�Щu�Րُk�n���{|��C `�85;*U��{:��������^oC�yu������L���nz R��.�����Dp��}��y�Ի��s柅��:J"q�J@�L X�h4s;g�����B�0�#uS3p����Cߦ_f�]L����U���5ޯc�֊Q������RחS�)gz/��<�%�rC�uW�@�67�_SnQ�	����� '���f� Mq�!���-�,�vje�1?J�\�) �{�RlT��J��}	%��[,��<O�P���CQ��R�k�S��_�yV�o��V��ndQ��}s��2��F4VCP`�X[>5}w��b.HNq�H�5;aZUE���uvƋ�J)���VS�ٿ�����#9tw� 1V�48(5��ʒ�k� ;�]x	��;~�2[�D=��p���Wt��V�!)��ÎX]���K/`4xee]	-��ޒB�X������}�☚��S6�%p�Eg;C�;��hڛ9D�^�]���[Y�u��G�&%���� �F"��KV�N�Շ�6����2�L��{���9��k�]۸@�eTJ���t4��X�5]����_�:�������#�[�u�5��u��|��b�l��S�,f����6}�1�y��k���"�OG⺭�����sD�	��U��	�e�GY=H��VK�KN!؊�e�`�/2���.mU�Ψ_|�Y�CO�"�����po�w�Y�9z+/�Y��	�u��%�6��W���:���=_6��K,"O>=�;?�%S�l��C�55wsס����V��0 ���T�k'Eaq��rb[ݗ+���"�X���ԩ�0R��� .�5���d�֏`���/@^�׽.���;��	�T5�w$�/Q�[v�����a<��������:ܪh������|{����{�{���Q�<��ʫm�>.�Su�ѐ�Z�����Bb�+")Bn
��t}�,$;S�F���<��-:C�~�1�i"����k4��{iJ3���#&�9M�Y?d"3EyF[k�.o*��K��4�ڹ�Mu~��=�}�G�'�|�#��Dd&��Q��1V%C+��!���kBp��w�ۮr�\��!:#A+�F��H��F�*���9f�cy������{9c�C�>�nj�l����6'��C��N_��;��*c�I��g�ʏ�So�����V��K�a����,����`��[0]mᏋ���a�*���;/k����j����S�'Ɯ��ҪՁ�c6�h�?}�4��P�?t�`�T�<��%��s;�G�稓�]�R.�u��HK�ew?A��WT���;) �x�_u?W"���q�IU�Cc�k�T�X�8�+��11��F&3�X�!��ɝQ�Ķг�*�I?�<�X�8���82]��g#�_~=~d3f`��Nϵ:����JU́7�4H�~4�9���~������ut�ѐ�)�_2{;�v/��TJp��ewoI��ބJ�IH�L䑥�wu�w�@O2bU�������f��4E�@�֮ڪ���iw%ü��8`��k1�
��"��/�825C�쌷�g�����]*����榭-�Դ�
�Mj����x�D��=�M8h��Yr51�%eD�:��k�OT�6S����ގ&�l}m����[�i����,}��IĈ�Z0˃Ǜ5�o�����!׵LԷ�::-���]�NXȫ
U5���y�ک`T��B�c�T����HL�2�"�Ø���(R��ؘ�*&ɘ����l��S�{m���tn��o�}�.?e�8Z~�S�ӝ��.gl�0�J	tl�k��F7bZ=O��v�2����E�u<1kr�4�݊u�Up�ţ����Hi:{2/gw��۽y���i�\�g���JH�+�Vk[Q���q�빼�ʶ\=F�c�Z�7s���?���;:��`�/�H���e}���8������fm���tm��'�I��?:���?C�l_ۉ.��~��#�7Y��^�|���f����

;Oz�k���>3�FO����
o(����Q�Q>H��Z�B.��5�Y5�xh��ړM?6q�9A[��A(�j��l��w�����!�u����E6y4�&�]p�r�u������8v7>:�&��]�&I�X�/���eU�͆�	��v��8}=�4��NY�jy��Qx	Q���=�b&C;D����2]���ã��w��s��	Ŷ�2��A<$�#"4|ʨTĀrlY�O�}K�nA���{g`���4Ҩlho�2�ĄoJI�Uݰ7�|}�]/��kր����t��`��cPW���|�����H�/��_��#979�4iQ�oB��
d���ج.����>y�C7���|�0?jq�b�C��f����^�WWΛ�)�-�M��$*�t��e��y�h�щ~�BF�GqZ�22J#�д��i1�%R�L$��-\;^�]�0Y�rw������D+�$y�� a�5u�x�J��'�̰"(�*��¯��?8�1� �s|1�#ZFb�3F'�WE\	��3%�b�nZ	34|�c�c���-o
?�3���6em��1���~r�8��ws�ğ���!�=fR���Fy7dUQۄV��jj���$��u!�]=��u���j�߳*d��,Wq�p
����?�)k9����3���P+VM+���yW
ʝ�ڟ���\&R?��Fg�xq=}P��A.�G�~Za@I�I��eF���w�9iAO][bZ�뫋�j6E���P�^}��Ԇ(��FWU2�	;�������Wx;��<�u08wT�&��[��9J�nK���qu��f��"�DT5n=bq��F|�{�ʎ����9[��������V�O�5�q(�h`�0<�s/���&��U{O&QUm���������?�C�=��P��ض|,�i)��B���r���n��;��)�sI�@�95��'�2�����V��o?���}C��˸z#����t��*#����EsEum*��-��Т�/�6},�Ф꾂�d,fw������z�=�oI*"��ZQ8�/W(��z�6���WZ��7�3A���9!*s^{|SH�Ɗ�6懾�P_+�����v�/��e�Ч�]��lm+�l���H��������sL~�ږ5��8k�ʧ���x�&��Ǵ;��j��%q�{S�z�}�^=ƈ�{��þ�v0$rK��>�`c]�d��=PpyRorIA�H"��xE�<{�8lmpaԘKZ1���Ò���7���!?��Xv�'�m��8�ra����]Ci�{�5���!xF��h���C�o�9�#����὾�&��SG~� ��]��o�<I!j�d��ƶ�27��5r��M�)��Վ�mw��U8Q��t�6�I��mo�hl���?,i���塢���: �53�>A�����UYХX��֞���[$�%��(%��Dptu���l_����`I�z]�������G%�װ���'���(�з�n�.��w@f^��M��J7O?��P+E�ͪ�ށ7������]U�{x����T�q50���?ߌ��7���R1 ��_�k�����u7��gg����w��u)�u�'������F<
�ɽ�^C+y���=���/�<7���3��'��G�"ޏh�mϘ�����3��� �]�ws�����`˗�%#���h�|��h���oH����&@(���E?��x��|)!��/�ힻu�Ƞ�k���`&�E�|ؔrT��s����Y'�{5�XP�����5�?��ٍE��[��P�-�z�\��z��"�;�OO'e��%Q@�x��G��q��	1������ ��vs��t�*��?�I=l����G��KUN���ѵq8x�1���ٻS�p�ue��d���Ǉ˴�Tb<0�-=:�ϥMy?u�LI9��rQ�]�S~qi�T�Oށk��c�����Z��6�k�w�]���^�t���t������]R�҂t7�#G��Rҥ��R�Q����h�6`�h��}���?��08�����+��\���\������HO��B!nU�T��f�b�^�,J�|�,�����y!R4�;��\��t�|Sb�gKK"ы�<�*��à���
S�Am��.��^tn	�	�}�x"~G%-;WP�T�B�60<;�(�ₑk�Ґ���C���+Q��`���o)�1�{Aj_ X~�p�^a��ѓfAt�N�=_�@"5va�j6""W1�g�hw�j�}�t?O�������������$�S2fw-.H�ԙ�f�e�)N��<`n�%��1��kl11�8����m�ȭu�Ģ��N�; j��i��J�I�	%�vR���P"�	�G#�;�Z��+���pڌB���6�{�$�d���O��
�<��q��-���D���, ߢ���ߩ�]_*D��o�L�7�eM��a��bce�~�ѡ;ڥ��i�u����-Fܖ���|�,<�ݴ��9���I�&����ڳ�(2�[`yr�Pե�#��:j���$wi/�1/�
�[��(���~�/dj1RY�S��W0��\ȧ����	��Ȗh���╺( h���`�_!��TO�c�&��\��=/�W��Ő��sct�[��`傴���˸LMO���U�Η�8)m+�[��p�s�@��k궷�9�-d���Dsr@�F&c�;}e�r{��<�H�os0;�q�K7�}e��W}�t7�͵�SW�P[�=i�64�ͭZ�.|qV[,Kɸ�Ɓ'��1�6�C����3�?61r=�p�v~���H�[=Vb|M�����B���P�U>şw����:=���)��xr��^Ѐi}M�u�L�L�P��R.E��s_X�on��*yK2a�r+��yە�6�~��OB[O>Fh����_�K-TH4Y�_��#�Jj�B�[ԭg������o�L�|�.���8���>����D�����W�B��x�0�1�r�}�p�d�>�L_�y)lgf���z������i�%.�H�@c��gR�x�8��c�L��ss�#���0�����e�^~���E�pK7��ԃ/�i�T{z�Ф߼19f�U����mG�?L�U%�E���4�L2���	$6��l(�p�QB�����{.�A�Q��ϖ�����&/���H4��^��8�;�b ��25F�7���׾`ߗ�W�pb�b�k�-��Ƥ��&q&`�Xk�Ky��2�����N���N'�S�,{�Un'|�q�o��S��I�/Kk��^m�R~�Ad.��wL���f�v݆��a��5�G��ľo�%�9�v��6M�"�i�A�e_�}��;K ��8�{_d��IO`�K��?O,����6�v�P�ЙYۙ���XY��īi<EFh�5K��FwG�gJ�G|���&3M���~P�[qW��g�g!�D�����uO*u�2�:|�_c���3�ٻ;3k-~;X��6l�C�5H$��#D��iwO�����.�
����:��~h���6N#� ���y:��$�����G㑛�d��d1Z�ۿ^�������ԓ@C�͆/�L>�\�0�^�@�D^�7�]��RM��R��2�Y����X2AV�o�(�:��߼!B3�zT'Mf�V�g�����lp�7},��m�U3��}o�EY�"�<�ɚ���0�D��b���43��q1v�
j�B���Ŋe�Y(.�:�ѧ��q���̌M�b!���~�f����������w�'��Q�����:|��� ��`�?n�&�OV�������T'��4��6��陥e�_`�Ӊb˷��ޗy�\dBs��%�]�1�4gb�-�Ğ�M���">�'2}ss�� - �#�R���F��sb�0�=L��4�pW��s�q���.�m�:�����)�3�_��u_��);�m�n�xL��N�WM�l��$A��֝4I]lH����$������%�1�-�"��3�})�h8��6����Y�^VP�nN��?���̫��%��u�#�K��F�@dt��1�=�.Ҋr���Y"<Tw���eK"6K���� &�]J<��_��&Dk��Jk.0nPc���4)�&�G��x]��գ��!�5�H��͠�(�nq���M�����`�v����r��+�8{*o��l���o���C��)�xy��s9�t�`�[���3��a���;>A���4n!�MQj���}8%>�M�`����b���f��*d-�Ւ��k{^�󌘏tn"�ڂ���:r2�3�����&�Ut1��0�����y�t;�/��'��m�k��@�V׈����=�F��fB�#ܣ˫p{��A�YAэ�|p�ո��3gBk� �
qAwg:ohȪ���B���knc����H����1^�{�]�z�c��x�����������iy&2z�ޗ�'�N]�6�l��~8V3h�S�S�?�n-�]:��Y_/.��U�Љӳ� 
�54	~�(}�����/�G`��[BB�Ĥ�e=�Nb�/I���&5�0��>��7��'"�W�l���f=q�L�	�R����+_��gBP:5���>��u�
�'�+��6���0!c��:�R!��{�v^R�C�%>Y��j�s�[.��?��3 `a52U�ͽ������C�2�#�n���9�Z�B>����~@���;���(bJ=7?(M���ɽ�gG��_����i���	��r#}Q��3�r?���	�� ;a�X��'�?�# ּo4r�)��C^i�'н�>hx�G��&o��w&�>)&3�0>r;Un09�&CT�d���;�A�y�j��de�����X�p25��� ��y�3�X(�zf�\\��Li��vW�,f�ɇ��"��	��;�I�!�>�(?{����h�n���7ί��_��&���R[��|i���^�:�:�Fz�yl�뷙��>�����+&t~�X��A�^��Z�,�1�,=uu!i����IC�PE�0ZR=;�a5�;�{Y�U9�Uu婭{{�� ��5��:$�Z���9眜���ۏ��ŝhɮ�\IV�g�K��(*)V�5�x�:J㕫͈����仟���K�N,'�\�1���t�GD�	'������t핳JA�e~Xk����Y(��?E\���i�<.?}u��a�i����#{1A]8""x�Z���!��4�Xv�����/�Y�E�t"���ڴ��FyӿL)�!�0����&��C>f�J�����
���~Q�c��FMͳ����#FӴ�kŹ��5p�W���k������~��n�zC����/� �m}@�H������+9@�bJtJ���C����4~���:�3��A���2Sӳ�`U���4�`�}���j���4�p�� �T��6'�o}~�_��
�?m��@�/&T���>�C~� &�Q�����p2RzΗ<��r�Ҹ�dT>;ӝ�w�d��S4��	k]�������^"�
��O�T��p������@�c21&Hij�`�O�C9���[��ɓU��w�֓�=���'�7�Y@pr�X�#�lf'ԽS����M��u'�V�Ե�>'r[8�a	�~��³����I���x��
,�{�w�h��QU�1���T��d�u���������rw��Z� knǤN^�j|1�+0�K������|���/t2r�k��q���v�e�#��o��M�ɣs�hV�c�8����Bơ��$���t�D`�|푡�v��/�3�_K�!��_��_������;������nM��
����+Ա-��!ܮ+���~�w�������Nl(�I�������j�o^&�h�Qj����ӟ�ڦ���E�/��ƑNCi/E���:��N���7�i�h2���M��������Ϯ}�U��}������B��-�ƺ;ᰕ]W� v�2u�q�n������l��p��f�#��:P0�}Q�D� �^}t�duN-��{j��R!
���`2)��"�?ow_u��-랿	����\�V_�j�Qv�����4z�5.���j��OqU�Z^�4�x~�ߨ���@e�7����E���汀��3�Y��&��Ny,NbF�i�^O/�%P�\v��i�����O���h*�����!6��0�h��,�3�Yf%��jhA�F>L�M\_�'g'�=��f8y$=���Vq�zM�0�X@�p)��������2@]u�"���lI��߲�I�ǰG�P�P�[�Ak����K����m]���z\k1���������V��V��}���g�r�l��O����p~�TJ�c�����R����
u���C �����Kxb��U��;�T�g��C���P�]��ü�x��+�rI��D�A�Ң�r��G+������;0j#%�R�d'\�^��ĕ��Žv�w\�i�m�Ǻܚ�N"�^τ�ȳ��1�o��v������XD&3x��:�S+*ذ��zD�:��r�䎓Yڊ��ҷQ\�ʛ֊&~�2�L\���<��8xlS:ʛ+[�L<ώ�(Tl�Ї?�#��231*��5�bf?<���̧��pw�s�����s��GS���w~,�n������uu�ș���39B��t
�['<����x�22�V�蠗m�����H�2�i+��Y�X�.��=P�	Q?�k\zay�47���կ�a(�X���z���+�'���_����4�:EfVA�[��	ғ¢��Do٧K��������C\2p�gh��?�`ݱ3��1܍-�ƵyM_1����.��-�-����բ��^��E���uD��ɿ������׏������v���"]r8�G�U�lI*W�2)L�w�Cj�w�r�.�
�,�]�V;�i�m��`^���S�(�#U���Ԅ\~������,S�E�5�QRI��*���cpٷ�8��օ�@+B�:ю�G�@��6
�91�w6�P�T��:�0s�-��~{�[��/�=ezx\�����)��苮�]��� ����zP��g�����b�^��׶��7���CN�h��?��kP���3�)
�m��7�י��_�0Z���{��,ʻ�~�4��o��9u^J9�Iʼ1e�b��=72�$�9#��@%��J�p��m�yQ.��p-͵�$���cU6DP�䴳�6!m	�/�P�p�Ѓ�!k]ｙK��+8b�P8\����q�as�l"1C�3�"����_w�J1;�O��r��[�2i����)"d�2ˏ��ù�d[C��X�N�*a̲gz�����!��`�|0c�R	
��E�H�BA��[�)����_��pW���i�i�G������7Z.n�p{����*�:VrmY��;Tß�p4� 2�"�w����x6�?2��V�R�l,/0m�mR5�c�A����bzZ�r��I� �5V��{d�zk�g�:&'�P9)EB����,�����m��s&vaH�Jo�y��x��1r�v}�˾IM�_`�oon����K��=�<㳫�lP5-��b������y�>JM���U�y�p�
�Nq=��t���}�b?�12BQ��K1�_�S�z`�䭾ė-
6{YD������DDFr9�<�����ۚ��2�3N[-�
��y��lp���z`���>��������&�q��}�"�oo���0	�F���!���K�hн<����a�f�yRH_�#g�R�y�ᗶ(�WI���ak"�Yj���U�̊���5l��xa}��sGq>Jih}�g��XZ�\��@��T�������8�2��4��G�O����w\����{�퉏�?���#��@`B�����EO���Fmˤ�������<͚�̺֚܆��_�fqI�D��X�:�:�����!�U��p3J@J�4���8=}ID����
��kp�@���]�]蚖P�iȵ���lk�� �l��5ؖß	�F)���О/�4��qQq{!���A F�7��NyU>s�������Q���[U�{���1��r��n.Sҝ>����_Tha�����x[���=�-�X����{�*�3�Q�t���_Z���I@���#�9��g\ɘ:�Nj6=	��z�$�� ��_��#�@B�l�­���ą#�U��=NZbݚ����d/��q�^J�G ��H�z�7n|p}]d������@q��T��8�%�g���3U%��a�����2�66��Α�!��
��k]��;G�5.Q�aIZ|-EM��Kv��$p�:/���cĂ�V�N�Ϲ��hO_�~͇ç��)3ۇ��[#�8�G�?��\x�ɥ�VFe����c_��̆�z)�>%�ft�+ƀw�*�pޚ����E\ѿ�c�!�̍�
�F�^��?��U f#ļ>7f�0�>���bL?�*�nt&]�m�/j����S����2�����L:��tv�Y�����R?>�娙Å�p���
���,V^r�\��:�0&ms[�o���0:"�~��]�DZ#�;F�?�>_s�����}c����@j���U�
H�5�,9���E	@K(࢖=<��'rW���������3Y����]���Z��Ci��s
��V���0�
>��3o�@AB.�̘0��zȭ�R�	U�Q,��?��)�����//`��D|b��r���q\ǡ4�`uz�%�rvM}J�C8J���!�I�/��H
N��"��VS\�,B��.�'��?`�������!J9���[���������2(>��=��*�û��On���nF��O���Ι�ǁ���t�<O�ǉ�v���8�'"���2n{�c]��?	�<�jq��/�A��k	���5.�B
tŭ <�}���x�[:G��.A�6n����7!ۆ��z&�+���(��m���_�s��nv���e饥 ?�S؏�-;W��*���	��ݑ-�o$A�t)�H^�Mr���3Ǆ��.����d
���\q��{�Y��~VH*w(QRH�̐3	Σ�R*Cz<�j�Z�PG6,t���5�����L�ۀ /9�̫� �f�F=���&ִ�}Ӹ���G�ZLr���qC���/JE���c����nw^�����J�s�g6�B^��ٽj�Y�=�Xe��߅�ͻ�n�d�>,�3	�
�
��2��o��]���<���q{鴕W]�豠`�?�ڕ��,!uҠ�LN9G�1ϡHnN�eJ�tw	F6�d�3C����m6������>��sE��*���͚	�9�E=���
�`�Zf)i���_ /1;]Z�l+����i�%�m��S2s4�ϙ Z�X���2u=����ъ����10߅�c�C��F����GF�?� KV�G��7zS�S:[����j��ǁ�ͥO��.������
cv�U^46��0#��)p����;Rud�d�/����f��Y}���5�����b\�x�L��*b�R R��������g!$f��A�?h=$G���^4��_<&�в��h�����h�T�3�M���?D��|�]\���`=�4�f���):B�B{c����st�1!b|�!���,α�KZoޞ�M�����7~�e2h�I�!�W�Z/�p��T6�Z�r�fػ��z�_'��uӶ\�_�[�R�B.��|	C�3�]ʚY�qN`��	)O�G�]s�qf�]F'r������.1&�@=Y��W֟���=]v�"�!1�?�m�^]��UG��oE�k3�ڔ�kQ��_��h�i��L&�d�+鱨�Y���qe���'f7}�k���I�	q0���]�����A��ߎӤY6��*�Id����ؠ���h��\3_A�{eJ��eUFh��<%j�+j���D⫑g�&��E����9����ӆ}g���(�7Dr]Xb���<棳�	��ԫ�Q���Je�%ÊW���+��8��CDL�i��6W{�l,�gm�Y���i3BW��8k��m�<��ql��qc�F�YV���${s�}���o#�M��0��h��N����9�܄�2�jV+��d� �s�]?��<��hzGH��z]^��3[�u\��Mu
rh���:��垟�p&����f�Л�i:�@`��Uz�B�W��W�*n���O��Ja��m�O�IF����P���>J����-��A8L�Z��ˣZ���VU��4�0�D���_�/'0DD�|��GO[b��.�Naf�L��!�{��%X��,>��	h���{��.�?�����,���w�8�� ��n�\��<�QB�J�/�{UX��c�YCGti��*����D��������X����y/��g����ĥ�g���Q]��:nR����nM���K�;+L��p]�,��qS���mt:��Թ�T�����|K���j`�Ĺ�aڿ��^�k�+� =�^^�C�-��������4���EK`�u��������F��������z�XF���k��,��=WA�����tgYS�sk����ے����"~�:��N$��~^x88�m�F=�|0<���Jv�/B�8~�3C��9_�rc�YՑ���W���l�^���\O�b���g(���4' �ө񋓹�����?��d$5���>.��o@ǉ�Ȳ���D���	�9��e�F����������4ۏ/���lC���sGV}�S�;|����ݣ
��)i!F�T��dKڃp\�4�:�H��c?�p֫�z��)��?@��{6��W3��^�jm�>w=���$�L՞S���Jۄj.	"�_Z�{S��U��R�����%2��Ap4w��|�B�s��Q1����ΪG��	m�y��r@草��b}���v��|Z�u��뵦�Y�b�r�M����%Kt������~E�ϝ��q�?t4	�Y�!Iñ8�Ė��[���(�l�<0��-�m����kU�N���<��7om����P�np�q���5��`Gn(�,s���J�ȁ),��o%�
�b鋈��a#r�o(��\��v�E��ņMw����(3��e�QԬ�q>`tft���&Ltln����A��|� ry���I�8�����+��"��X�� TT_�G�d�tW1���D��X=M'����}����}����Z��x=OՀ6|@�XޕT,Y�XX�O@!m7~xS'���5��A���/��*��w3-�'T\��V�_t����P�+�=+~Z���S�K��ٌ�c���e5�G��(y��U�-2�'[#,��zC�8���^��Y��l�wH.p�K&�p=�Wh�����MD�6��Ɩ���{T�Vf��%M�U��Y���a�W9ɩ��(�l����j�BDP܀.��8{�_��tHp��v����v��0�I��қm�h5�M�Y��1���x���oX#�cH_ϛ�Š�b\�jc���8c� �⍉e_�Ǎ�������S�V�n��]Ϻ��sw��h�Q
�+t�U�l����6��m�bզV=����������

�C����8����v ���\g�\�R|��
�F���{��N�����I��Xű�Y5�hy�/V9=���:"9�m�)�:��U�j6�l;_ _z5v� ��^��jn� ~��#��i� Y������QfIp�5�@��$`�䢷�I�JT�(]��?�`�Z���������re�I"a#���)���*�:Z:_��E>Ǣ��w��:w2\X�	���m���0����&c���*۸v�l럻����	_��>��}}߇���e�կ��:��҆[Z�=B���؀u��`kD��Y�0�Dݑ�5N���k`qt�g�e���r�N��M� 1(�W���Z�|�#>0�fV���1�@UG�C�>�1����llG���-ty�u��gٻ��Ա������՗�I����}����n�����v�]���2�p޵8�;�a��tڏ�嘸�Fx7�C"�D�nμ���8iMd���eL���9��Y�k��Y�U�S��(����cƟ�2q:O�h&f6�ӂ~h����!�-�]ؖFF���᳡��ùSj".k��_-�Ɲ-����\�U�G�:E�Ĩ�߸����������<
�gb�Y)�Π?��OMR?"�\�	�2F���1wf[�}����8&@��Y�&9�>U�&��]h��/�ɿ�5�+�-��㩜�B�v�c�7D8O����o��d��5���bѓ��{��\Z7^�ڻI��n��P*�is��8�p_4A.����j-ϼ�N����hb2��~h=^YШ���P�ȺV�W'3��Fbu�o��9��\�N5 ����t��i}|+ =:������w~p�s���PM>(m�Q��@0����c�+#aۿ���S�w߲�w���"������N��v�/��ܗ��=�zB��!���,*X�!0�O��П�΍�X.zMϘ�G����,M~��=�nѲ��|!�nא�:��O4�6�잢%X2Km�!|(x_@mk�
��B;]_O�e$m3���L�y0B;��������j��Ɂ���k��Cb�D�#�P��2�N���l��i�ZZh���~�d#��Ϭ�N�}{�}��������hT�|w����;���a�,UD�m"������ޛ�;�̾�tߪ8�>�b�����htϩa�bp��b'=h-sE���ţ����΃�)�s����V�Hu�Ꮵ�˽3ȥžl}aG\��"��++_M���-ҧ�xdL��H1��=d�Ә��X��|p��F�g7P���X���b�@D���n���&՘G]�iJ{�Ko�6J�O�p���a��#��=ضF7F�;�t�}`��M���m��T�0B����ɻ���rEÓ7��h� �\��G�ȋ�[���ގUN��Nπ$�*�����*�bp%��'N�a�������(�3��k;���-�b���Y|ڃ�{���b"tf�k�=\��ʾ�nLP�
D���
�K���Ţ�'��>,1s�~��+�A^�d��^�heK.��Hk��q����J��"���C��_5�^<�$�W��ޙ��~>#yx�|8�ȹ{��W��_�7��O�2h�K�����I.�x�_�@]tϻ��b �Ɂ�`6�=ˍ^���/�P%�	���l��_���c2�f�z��� u��BEWU
�l2˝�=5��X'hd�3R¼H�;�������A(���n��DZ���]K��Ӭc�ri��3������Q�� ��&�%]�7��
��D��+F'ߺ_�C줣�!��;�a�ՠ�W��AOCL*��Wu�!�hA��w�~	[��]�Wn;,|;�~v��6Bu�s�Dy��n�����u!��re{)Bb�x�e�Љ��|�(��X J��L����B�Vx�`�9\�Z��W�L}��n
�� WW��};�v��������SX�+�G�n���G�U�q�cN�W���k��b��z��O��z�b-��x�6�e�7��:�J����eꛞU���¡�q��<�3�Z��O;�v����Ӣ�s��� N�4��'a�}ɍ�l�`�an��9�l���{-|��;�33'�it#��ר���N��:��7���v�㒌o5�]�{UQ�EK?��ncե��s�=�@_�z�/�A]�ǹi�k▘��+7_'���N4���
��b�^&ŭ {)~?�q!M�A{�����L��?4�F�ۆ>��L�	Z n��i�2�)��qՎ����#z��	���(��ܨwKC�8Y�T+������h9��|��he�G��L1�
?x���}q46r'�=�`��B|�!\)��oh-q`�̝��ж�����"U�1����~�DxY9pP^'����P(�-�I,�����x����G^D�իմ�z&�Z�q ��J;jA�9�B�SU�b�KYI���g���{sH��h���C����/��_N�%��<Λ�Tú;�/��_�=�g�	��P�Jqѣ����a� G���ݧ���� ��>���n�7?�2g�R�1�4�i%U�eo��X��~8��Kn9�
9�3by�Ԕ�J����*��7甥@�tBD�;�����.oF�}v&%���;&�?f���֏�ܘ���}�q�^8�#����"��':�0��V��~��J,5)_>ӎ�&/�?-��ԟR.�dU?`��8a�	a�_զp���N	���{��_.�і�,"i���*
� �������Hw�̔�j��t�1g���]C�ݖ:	�����T�$��Y>7������+da>�,J����`.{�0���Ժ�s���r>y��v��N#�3����Q����ɩ����X��F����O�V׍������a�4�4\+	
�%�ш�����\�7N�%�b�?oH�;bL��5����+5h�T�/^^j�*���>�8?}�����(
��v�.Q(�G���WAi�.���?�5u��ޅʅ�g�4��h�o��1������{�����o��G���~KG*A�ܪ/g�n�+��hL}O󍵜S	{�J<Ck'��R[f|��'������^�\w�l ˽�NN ��]oah^��������=8+�����>9d�|TT�t['�����.�;�t8�vGp;�5�އH����8��������RR����i��67��J����9�@4F
�F��p��;� �tXFv��Xi�(*q�+�s7z��L��|��HA!�Վ��.j�Hh�v�Q`���~ �1��KL�w�G�(1�cGi�KfV��2��L��LhJ�����G�C��e����A$p��Uf��H��5�M�f%3�pQZ����g����z4���eLmQr 1�o��3�c)���R��`���&m�����/��X�{�qA��S�7�>O�9��p�@#����ֈ����I����Y��w~�ځ�U�X��ʹ����� �FبQ����QgX�^��1�{���	�I���EC~)�bÃ�a|�Q�,��'r���<�m�3-Sկߺ�"��8�o�V�j�.�ON�Q���]Q�<��M��G�*�T�g�0�S����Rt	��6����Lk;S�P;2@�3�9��Y�Fu��?ʂ��{V���Vu���[��'(��~���v#W��.��`�mu���ת���l�[i���"��;����+���~H�]�zZ��t���OI�o&V��!�餒ള�S��a�R��I��rL�j\VUqx�����G�0|��r�����P2�2pN���o�����3#P�"�������I�������B�d�3�n�xW�v�I~��CCM�����9*h�ܰ��O�z�"�i�4��(��a����g�S�P3�^����ƔԢm�o����Ы�lbX8������Dc?�C>d�2�V ��;	{�<	AvU}��FW;C����>O���;�7�a��A�T/~��v����^��]9v�r�|/\�����s��nZՎ�K�'�h��9\G��e.s�t��А���K8�`Yz	�2��J0̈�u�p��L�*�M�����rt�S�ǎ�׿m�wT�����M+nK�����U�����a��h|<���<EU�92�������9u��Ă��}����j�ȧ��s��	N�F�?�e�W����i
�y�M��K�����,�KNCw}�����5��X ��Yr�IW,��_��")[����%���l@�V�t.-�?��#���z�OD0��H�!��[d�����g�u�g���H�y���,�!,\̹�0H�U�NO�{RS�:�e�j�	},B�ʩ�7�*?-�s?��]m��|3�s|���.��ˈoO�	y��TR�ޞ�_f��'V"N�Dh��f��?���W�⪱�=����)7������:Q�r�H��\��#aXP��Yd�Æ�P�*㢲�w<?a�E_�_�������wu���P��A��qhhg�۫y7ٷ�K1���[�m=L�B��<�Y�,��#��ܠ~)�/Q@�2�P��G�p<���0}^����L��
"��m��L,Z�϶ɍ�:����kI��W5%Z6�;�V0�&!3w֞��űV6p_�4F��*�������\@�-�]���U�:�g��U]�G�٪}�]�\?�6ɘ0�h@[���KK�U�.tv�e^CY�4а<��<���v:\�E�v�cO�`��UT�󊦒�I'��%|-���dl��.�A�Κ����@��K�Q4�S�UB�@���\��	<
#i!��H�,�&���A��~4�~d�ueU  ���B}k�*xř'�n�wF�H��[}��HUE���lc��W緎)�i�˳������1�}���" V%pQ~X�k�|�ŭ��+r�?r�h��J"���-��bZ���9a���N�\wt�=��?��;3�̸h2�E���P2t͇��O
��Qc�b~��v��v3~�ޞ(��>Z��[δ�94d���L'U���wE�k�����}lE��N-ð�`�Q�M �����	����%���M���V��XO*O1�W���K�R �]�Xn���kQ��p�}�cB�3���o����^��	�-�	7���K�k���_��Ep�̈˯��:L��_Z�¤p=d�ϕ�Gi!v�9q�Ż;6%Hx÷��13:TqX�V���儎.��?�O�X+7��u�E��-}�v]�sjp��֣���8��������]੗斦*<����D���o�'?v����^�Umt�\�rWl���I��%S;�L���6h�Ql��rQ�1�ڣZx�]�FK!Q=M��&R�\E��W�O�f���
p ��.ޜ?�q�1@�ݓY���Y����-��{F��뷑�����K�(%E�cY
�Y0��Q��ޫ�+���\������,2��s�~3c����ibc��G��l5�Y��vڽe]YD���z�k��X����2��×Nt�w#��Q	E8.���1w�M�?�=��bϹ��M��7t��8|+(vn�:����O�@�B���
&q�!�3�;�#��ƴ"�jx�&�r�>u��ǁ.�Һ�a�Ԟ��^@��FU)��V�n�����'��L����=)�/$=+��N��H!q�8��Q)r8U�+��fb�uamU}�<W�wS�>�8�]"u�뼢X�1
8�JJ�ߠ#�
i�&�V�ۮ�ȍ�zb��~�f/�O8娴>2����1	�9�)���S�������t\:{�h髸��d��6����0����0�ы��i}0Ҁ�ӈ��'m����װ��;,nԅEj �@xV��J��I���';�L�a�Ef�<��^��wć�؈�(X� s�;d�u��CT���:�/nz	�c�&�ٰ��[�Dv����X�D"���bzp3z���& -xVӫ����D����Q�e�}M�����'�i�eI�y��޶a��g�]��botZ��G�n�&ںdY=ܔi������c �0�h� ����w#/�I6�,�Cƿ�Պ�2����H���l�\jý㇞��԰��=�͖!��K�طތ���~������x����vԀӼFX�R8?k�����ˇ0[	ϔ"tӾx�)�B��wg�6a�ލ�����۱w��8z��	��;i <h��?u>^�Іic�Y0��� �N��-��5��qs�~�z���X��zY?��)�SS��D����A�y�MH+�����Hڗ����C�}N�����81:��N��у�!t���>�P~'�dE+M!�2śd��v}aQE�	#"�	��X���2�C���<ٲ��e���S3�&������V5�l�+K���aaF[��oq�ADt���7{��c��q׵j�cڠyyFh������	|�}o���rD�1���r�4b�=S��B��x�{�f�j�	�	�
�
���ss���â!<�惺�w#2~1�D�#�Z��#m���U�E�:�p�C2�L8��*]斑 ��v��9͞�'J�<���w�@4�:���&U����ބ]<��K�k>������W��*����N�Qs1 uw�*�TX��pO����,�.��
��&��6�91XL��CG�\�$<��s#�	�=�1�eYgQ�u<�w�ks�A�k��cl��/��O9Τ@��k���t�6
�s��� �(ͳ<�-�r��+3?�������x饒��tT��Ղ@f�G��TƔ;㩆���9_YE�-��a�� ��א.��ˏ�m[`�'�]���x�A��(H��z@m��J+
�(�9��e�0��B{Y����i��n�����szFj*�v���|jb���LF�K	��Ś����o���-�L�Z�>�ن�li;)D��jg|�L�,$���n���!���i
��d]h��+��~X^�2�������O�0m{���]4H�d�N�;���xDe\�7�Sڕ���eV�b~��	�������@ĦN .,gUh���xu�[_��\�jYr|	VWy�w}�_ڑk=���J�<�w8����oT�5JkV�"Z{�a�5k��;�)UTQ{S�WP[l���-�g��b������\�/�u�y�s���y��s�E��n�s@t��L��y'�:[('�3ŀ 4Bq11C�����ů���AX.��
ą���v��;fn����*���.3v?�eq���L�S]�Z4DEcBN�^��N�xkt�Z�����Is���͂_/�l�n�=�8��9�r���߉�p�>j� صS]K���1�l^MY�N�tW����0�r<
�\$�^ $s9.��O���͵����MxՕǧ�=�\ɾ��>95vB3�o���������l~�f６���M�J�x���ii�ƀa{wr}�[hċ7��}�,�˙<���NQ'�^p��X�Kk�GYƲ���/ֻ�=F8tF�}��_e�\���(=�o���'���ĕ�<NV���[���P˯� ��&��AD�F����j����(5�v�Ζ鬜��@7
��~�1:(8n���˸��2�y��̎�_+9���2L7Gq9ܔB�݋��J��~4]M �����w�E���A�l5M�|��DҶ=Q�(���ޣR뾝V�N�Y��/g�Ǔ5�QuL�ԯ���)W���?�bU�4b��fP�'�a$�.����v9-�p抢j�^l4T�:�a
��d#ڱj�z�D'�E5��3�����dBJJ�12���*���T!B��T��on�k���"�j�׎ߜ��-�ch@;uy��������hq�chP�g�M�X���a�%o]'U�"	l�S�m�r���^��<΃Fѹ��~q�+}A��\�P���!t�k��]�H��h)`�I58��x���xaW�zz�α����r��f���ϸ�٩�LV�1b�j���^t� �8���~c����h8��8:>�W����үsDG�݅�U5� �J���/1���c�k^l��) �#!	���=C\���+wH��ɳ�8��9���0�/����E!)I�x����Awː��<��>��߆��lE��a���B��D�FX=��3���TĽ�����h�5�%0�̝{|��_F��(���S�9<$zhnnD乨,:���C�1�����Df�Vp[P(���~�����z���֚�\fr��ҟ!@~q�-Y��1�UfR�Y5f C�����A�����E9�_���[K`4�Y�p`���B�);s،`��z^�j:�{�L��lE�7Ʊ �xSg�l{���OQY[��x�~x�i���ћ^
0��·r�E[��K±,���}Hn3b��f����PN��`���B/O�37u�/�V�[M�f�v@���L?�Ѿe7ԄFf�̩��Ϋ	9��N�2L�d&�JJ����� @�V�z��|S$b9��>
�:�
�#_����J�޲����m�'/%r���Ɵ��
�sݚ��sW�������߮�S}КM�0���;����s��D������#���=�k�-��!s��@��p��-x��N=��$���I1Uܰ���^�E�������Q	���A�	Ԝ�ő�t�H䚦	�Ea(:���\�� !eip`$"7�)Us,C0X���H��J�ࡓ	�{E`�N�~��}�W9����JO�UF]�:;��8Z^�����'�tᗪK�`�3����1Bj��<NI��f��MW�<ֽ]��W�9��)��m�_�����Օ�^��-N��/�t�����A��2Eě܎ʲbN��>yY���1M�PvM�j5ғڼ9���6�a	
u��75y ��	�r<�bޅ��_�ޒ�A�_�u�Iz���ZL��(��CԱ�����{�;J޷ME#����P�A���\5rr���d�s+��T���.���뛽��".S��:�߿���L��"�,=`.?3��1i�Ao#�2���^9����f_�ߡ��\� `���'cͷ��a`��s�׮P����y�V[x�cp*�� �����!��W҃�G�'����D�I��hEK��M���*��&,%�n?���YS��}M܈�3����jʬJ�����t�mh�e��H;��w�c� ��8�'j9_+=|���+���+��2����X�j\�b�e���G����߭�v&C����B��YD�R��^����S�l"'?O���>�Y�(�Y�ـ��[�M�Ժ��3`��q���7�ê������T�����e�&����%�~i�j�`??�I��� C�(e��m�Hy�EX���h��C�1v�M����؈�����c�'�A5�j�7{f��#�f8q���D��ڠ�-֣��6p��BBf;jC����R=]]��O�Ξذ <o!�Qt���Ly3���gj��j�R�M��h����ϥފۋ�/�&�{�Tg-<����g,�)��.�c���4E�6x�U�d��N��T��g�T4I���n"^2�����I)�}�1؊��#�餔$~�.����$W��N|��&���U*]o������c�����XWpj�]�
���$?�-Gg{3�5�{���C���f����)���=�����-G&XP\�Ҕ%���9�l�{������j���>~�u�=w�C|ˉ�����))��g,oDa����ת}�m��S�Z��X����"ES|L)�9�ݠ��μ���+��E3�����[��F���SE�6
���ƛ�ޭ��BF}'B��I���e���<q��ߍ��?��3'��w�:��D�Cu�T��J�Ʉ��(M���m0T8�-$�1Y���_$�|w���2���S��67�(��UJ��<o�g�i��
�t<N�^
�k��Z�.{��eI�V��O�*�)�Q�_x+�u�G\L6���+
D�I%�p�D�	-�Q�~��?y�{�|��(��S����}�"K����ss�r�}2��2����\�ܒ@�- 4����w_��{77��>�oh
�������~REE~���}��|�J�p�1q�@�ͻ��7w�B������:��V�N�Ka`O����cnX�堤���� j����&����o���Y�~O��)�=v��1[�*/i4!M�b�^���>�la���	76��	L�.O����O�m�@����x&���L}���y��}ʰ��T? ��:�>����k�z��a���VR�=H�`#Q�$�flw�[gA�t��L[�u}u�|��{�V�������-L�;"�<��uc0��+��VL�b�F��\{C�\���Ht�U,�������{���ϑ�	��M�a�/םUt�����fM��N��$2sO^��V""y��t]��2fxC]����� ��D.��k���85 ������;�^��n��c���j�1j-{s�l��N)�����g����A�ų��k�Y&���6�*��d*��u��:��tA|�"Y� {�%BN��l����z�44
��Q���J���OtJ5���8��cy�VH&X�l�V�>�qt�
o�z
J�9�8[���ӅH��H��n�I�n!Q��ʘ>A
p�ʍ芌H��d��b�#<�:.�Ye
Bѥ���e��]���L�\�Y�Ch��SMQ����
"�ڛ�$+���\_ߖ�TF�i��k��_�AL�g)d%b�b'��t}�g�9D8dMmβ����7�/�d����8�R8�q���l[w��a!�������4�>Q�mcnX�.;�htm�gY�����Rw�}�4)a�<��{�]�Ox$��4\$d������9SIhI��ٖI�D���~!��0�NYn���.���z�+ڪ#`��O�}ȱ�`�'��CB'^�joi($��f��{j�w������U��L� S��w�Q~_Y̿G��(�#kvS�l�R�XG�8�!F�gQ����k�%�J�R��xL�(i�4���t�]{�-q���.!)m�����Nh�+�fkoZ�#�>5��b�N �W�_f��n_��8�P�x���&9g;z��hp�B�.Q�ͽ�İu
�����o��X�� ��<lL���m/1��bZ�Z��-��M�?���8�Q�݇ ����XW�<�{�;[�GH��qVq�D�����߼Z{H�W*-���IzERO����?x=��AS��^dA1���+�
;�m��Qa�E��$h[>����ż9���,q����uhO*�����̔�75t�ɑ��0�-�⡾׷���'i��o�OS�)i�ee?��wvY�����c��*�q}���*�rh�T���l۸�f4���$��<���A��h˚%!�#��U$7�Ͽ�ۢO�����	`Do&����U饅�ǅ�l2긘%:�k���"���;��D������(�
q��z(R�������!l2�3�{�P�
��*��*̩�R�J�����=���P��r�� �=�A��^��dl̤�N	 K���6F6	
Iw��i쟖�-���t�uI�,��/����	�8~'�ι[�+��\�F������o�i<��b��C��J���xBډ���?�xYE�쐝��z2P�+�~r_fE	�;���s�q1NU�.wp�2�����s��*�/���G�����7{�8Ga��ʹ����!?���k��KH����@����&_��Ɔ<N�?���#S,�O��3�I,yh����=�U���F���c�2�����b��3���%�4;;;W�T&V�	��_Q|4傕�1��t���S֞0u�>�-���ݤ'�(�o��x^AÖ������[~�|�����k7��B2a&�i0��?�]�3 j?}&�X�>ܼA\�����ĞM��t����T_���X����`$����O���]����/�� z�M��}e��L pV�L��3�
��U�؅��\�_�\��-�;����bϸ@���K����ۼ'��Լ�.����1$S��$j��̏R��_w�5_(EȝH&���1ay�$�a�&k�8hVA[eq����1C�z2!c�3��(���5+K�Z������&��]�J7�Y� ��+&Sc�1��˻y�������Qh?�{�z�g��.9l,xn��
�Ͱ�k����К��8k0�i ��ᶴj������>�h��v˄��"Y[5��_zV�ܗ�����.��MMf�u>���:��Bw�z�KqP��U�Q?��'�\?�9Q�Cȴ1��@�c0�c}5k��4�6��*�s]�h]���0�ZQYj����
����)�w�Ge75���1�)a���979ƭ`��V:���Z��65�M��&��� 2&H�{��؉�o6��{*�$�
E���,P��	���%N'*�9�U�b�߆�f!+���\<�h��߸JK_nޜTmਊ��Z�V�8u�Wzk��gϋ��/�P����ͣ�ԏ����
 �G]e��/$P���8�!q|�����Kg�}�|R�kݫ�U�I�j��=?=��_yR_=�	(��<5�O�߇L�U5�I�л^լ���=y�ظ� �-����Bh�qv�gA(�H!��4�?�	��~�Ul��o��~���9W����ÒA��IPd�P��5c�ca����=�:C�a���:a�ϨtCv��%��l��>����t�Ff�e�d�]�ڙ2�@/�<�G�^K=ґ̀Y*����N��q�¿..��N�ݛ��?-QM�2u����M�o���Ñ�'%>�1�P�ao�(�����.�P�����jW]M)k����n�^8�3���۸E��5�w�v;���t�"-��ۤ߫����a	oyvÚ�pB2�]s��2�f��9���C��� �[,��A��%�A^�Fox���?p�`R0�3~�y���a6���E�d�m��`s����ʾ�㥅�Gܧ����J�'�Ë�#�ݸ\������EQ�� ��N���w��8���ٞ1/{�D��<�_�X6���g!��!y��Y�qf��5ߞ4%�x	�1�
�KZ�2�;nr�;�}c�r~����dT�	I����>8�Tk1��@�������o���E�4��Օ��+�ᢗ��"�����T�]ŗ�4���:x0}qǩR�^|s�!�K��^�T2�~`]
�%����7�l�"E�Գ�X��>?��Q���`>�;�?q9����qW��ڗ�ȼ(�MR:������f��R���E�x���9tl�Ϳ�K���l��~FR�4�CW�3�NRwO}��#�ܾ-v��
�e^|���=4��j����J&ݕ�3�H Z�T��$et[�	X\�e�a0�9�	Lyn����.v��yO���%�	���<��+���Et#��9��R
r6|���4���˵D�6uS�1��F�l�ֽ���"��Ԙ�~��<δ��Ο���ԭ������L�v�l\U�2�Go���]18��?`;�b{��P{{�'�s9�#��d�8�])��F]�ߏ�G�K��n��~@Q������S��M�'k?:����@pT7f2:h08�����rۖ1�<L0	V��S��	!+q���2�>9y�n�N�oa�|���j�zGӑ�[z�aI��!\SDWk���S�
4eܰ\�L���{���;����#�AX���Z%��>�g��=���܉G�+�oH����WW�$�E}��y�,�I�\jg�"uI�X�4Y�1��+�ؙ����~!�'�ѦZ��>X��;�܋�{�ɻdl[�2.�_���qV"�䲌M��6T�"���|e� ��U5����K�?&�蠵�mw�2��7n+�
�3�8.(e���X)�s�B��6�OK�%z%�4g�S�<ꁮ�;Qʏ6KX*�����]=��v.�B;S-���e0S�p`+�S�@ǒ�t�9��lVx��S�T�L�_�wǴ�p����[__}B�KZ�7�^s��a���j/�:�K��C�lR��j
c�#����O�td�sk�׶�_���m�!�)*4�<������3����`�~[=+{��ڏ���H��V��n+,n�o�>�P�p��z[ɕ���h)tx��{_�4�r���*�w$VZQ��w�H��k�*�h<�:ۢ��Be�Ka�g��Wɘ��$�O��|���l�*!�a��Z��ʱ��c�k��(��a��OS��[�����Ic(>�>�,��H�/�}.�EVv�U_�k�h
���A��4'h&�W�������c"�ap���G�$�/������h�R���|�V���a~��
��&���T6��+������,� �Ul$$kj@�P?g%)=q�i m���){��Y����t�t����*iMd���Z��J���Q&]��{A�fO�AH��(
:e]��jU�⡗�����?X����4�~������в�Z[]��2R��3���}v�6�@cQ �DK�����1�{���_z�8�b e��t��n�[���&�2��=>�� ��ѵT6稔�Q��r?|8��kL��n��Kt46"�
��_�=����2������WA��Wh��a��v4L�Ƀ|l�?כ6��[�.�>y�ݥ�NRFVeV���g�f�U�)lh��R�#�#S��m��('��#��A�r-I��d�g`Q�Q����{؂>���h�V��d^r����}����;\��h0_\��2�aX{��.@��y�犍����;|?��)���]#�9CK���������|3�tυ2-C�e�kw�]��3����� R��#̥�u�Z�[�v��i����q؝ �����̏��	.(N����>�}��T�����Ӏ�>1�h,MܨK�'�Š����	/��o��[[O�jQ�Dէ1HҊ�Š���O ���?��0R��su�e�E�O-����	d .�oW�1,�e��j)�6�]sc_�1V}kl���Y�m�ʭ�hcO�Y�eȎ���a����L�ppT�3NǦ���֫%F?:a����ԏ��%.�{��(C�I3��&W�|�V=:�'ϗ�5��[w���i�����8HBr�����@'Ht�H�hX7�x�q�Oݢ����]I�x3ho���B���S�[Z��o��{pƉ]?YN�|i��|\�8:
1�y���`�l�'��I��Z����K�&���\C-�-{�T��Wյ��}�u�u�+9����1A��thj����n�z�x��6'�{%Yo�5@E�gZ?j�M�����e�O��Q�4�_ʋD������^0ed��ZP���n�9���F���(B���\`s;Z�%ͅ�2@�͏p�1RM/�Kʭ�_~|Io~�����#_O�^���3,z�'�܁4I	�����n�pp��6&z�}��a(��Į+-�4Z~�\�9�ڬ���j�W ^�'����6x�����UT��}�)�J9���'��Z&!�R�hʌ�>
��C�-Fc\dR�r*�P>P�Ā��k�*�hG�\t�j���fT��;j濲��3����S0O@��l׬h�4ɘ���� ������]�� �f��si�K{��g��5�K�53e�}ó+<K ��v��V�r������UXkxMwOL_P�*����lB�[�4�tJ��;^@b��1>N�-�Ԡڸ�}UXZ���ͷ�p�>)��sz�=�ŷO�^\��t��ߞ�}������mê�cv��c��H@}�;�L+(Cx�o�ω�G���Fx�/�Hߏ�X��!�L��`,��S{`$x�!l  �1�4���a���O���k{�"C���+麆2:#�b�4��u��[�"R��^�&�w4�7g=�ú�V�����L�\�e&9�6S���K���C�qimh5�e��@��`������lS
�~����#��X!BA�+Ӹ�J� �o�\���~�߿v�h�}D(�r�4	}1�,8	��m�,y�sj��6����|��!���噙��2�_t֥��AA�`�|�d�;7��yH!�-+3v�'�v~�G��68l���%S*�_&�T�
����N&�ا#��%�{�e�u=m�DHT_��y�5T���/��W5��$������\�e�ͶF�^'�R����ݨˊ�M��)W��'q(�p�b�Ϛj��(�:�Ǝ���֪�sF��9���/���=g_C��uL�	k��e���]z�#�I�����4��B)����Y�n��G�`2)h	�f`��!e��2^1;R"j@8[9{#[�t�3�%��j񐝧� ��  ݚ��Ӈt����az��z�l��2W���˞�"���b����>[��]�@���lb���׌�	ppX#..yᢳ;���=�%��;%ξ�+�ʂ�k�ˏ�"���^�pp�v0�ˏ���9�]L
1G��H�hүw�.�4me�f�;JQ��N�����6�ơ�]&�T��}A8����5�k���*��M��ee�W�c�:�'��+yY����^���i��~�;}y��MJ7s�޺b�<���#E�6C�H�UZ���|q���Q���㦅��&��d5��>�"w�R�S����*�hKt��(�����N�� ,s��4�;I1��^q{KcC\�96���%�}�4��I���|e;dW�>6���i/�<�U�89+_����n��=�z`~���mni���ș�?��;rW�c2<�����pRMAL��(�u�6ǿ���tO��Zq7<�� �f͒6ђBh��,���g��
���S+"�tq:��Y}�*�'�ͦ�?���̀��JB����gl+�߯�"�:���Ƶ�oP/���m��A%:��W��i=�ָ���FW0������,X���VQ)Q�ES��L����lJ�z���+�~��v��������d�eТ��D�q����~^������m���Ӏg�Q6
��ru^D�s �R_Xכ���.����}�et~?�9��Z��b�Z5�TR����]�&�=7V�I��[t�$���n5���G*s����E��J�ݲV������[��xӨ�}����t|A�9TOq�G2θ�>�V��E1���_���������gG��z�;�ݧ��ǜ"?a�.�7-�õ���R���~O9J��4ڤ��H�&WRW�[2b�"��0ф��mn������>k+�ML�^���]�	O(6�����Y��� �'<����;Qj��ߢ�]c�m�{;���$:����m��]	3���z^1����G�8���<�p8��p8�-�8�(�4ez�V��"��^m��$�+�m����]�y��Ś�9�L�9z���)1��6`�4���.�K�/�$���<��3���672�sV�!�Э��%�%���o��:���o"����3fך;
�����Y`Ҭ��g���� [�s������u�x"�y��N@��6]Tv�p��&vuQ=�~Ta�5�jx�LC�'�;�����fa�����N���u	0E��ˑJG'ž�O�]���!p��o<j�$%�d;�J�{�b���TpHg�t�a96|��0-PG6c1� O��{�_��a���\I��F��Z����Ʊ3?:�����b���O�Xy�U����K�4�e����^�bFH�	{�t��5{�����QpN����l�Պњ\'�A?}��#Y��5'6gl�b�=+��c
r6-���;9�P66gj�O��3�:pg,)���8������B�4�8�΃��r"A^ ^S}v�C�#,s����tM��'���u���*7����H�f�z4�,�-�����z]��ggK��TEK,�ˊ_*!�X�Z1Rqy6�s�Y�)}*R����v��|2vTD��ظ�5oH�� T���Z�+��;60��n<(	��C�&�^ش�|���A?��ao���V��?�Jsw�2�$���x��3�������`���f���6бLj�b��߿u��7)����YZZ��H[SW"����F�Z�??���5��6+Ȍ�!��`3e=`��L������]�[���K��w��pI7��������Kx�EÏz8vF�,��AZT����d��v(��1��՘Jۖ�#�����m٘����Q����j�g߁���j\�v<t07.r�(?�=��R�g�R��ͮ�Q]ӿ7]ù�U� D�m�wB��ѻl�t��(%S:jg
r
���"W3�ѝ�6���)3Z�@��_��|k?�~vh�gM�TE���M&���a;�H;�|�V�����=v�s�7[�UN��d�4��E��H��ܷ�^	x_�722|H�S$4<v5}v!g��)���f>ݯn��EN,�¸ ���7g5Ɵ2LEe�'gLxݴDJ���VO'�w��XR��{;��y@s{n��Avݠ7��p�Eu�^�t�Q��=0��9��aHJmA��wŷ�k;5��`i�y��b.bS݅Ӥ��88�X�p�}�uT+�k���Y���=f�42u��a"������1a�9��C�7}���zu#��ĕ����7x�,/�[�Z���)���#�"\L�pGH6R/0��p��'.���E9ǐM���lSٰemѬ=^��2S"�&2�8K�(�Z���{˻جZ��)Ԋ>ld�^t�Ӓ�0�s���f�F�؂���^-���^�J��2�����l�s�$�'��E��"��4;�Ǿ��>(��Uz��~!�_맋��X)����l���Ϸ{m2�����S�ً���R���j���'��Jx��r�d9��A+�v_iY���Q����a11�F�(�Hqe�7&�ox'g�&�������J�9f�e6���|�H������$J5���dD��o�qt,�	�q�]v��)�Y�+<�C��tU�%~�[��>���a��	�>�_�O�I�/�~Q����gPqCF�."��G��.���K�G������[����N�KR߯O�_�!T��
��R��\}r���Z�<�z�%��
eهZl*>��ܲ*QJ^��}L�}������Pptє��5�56h8���M�v-K�p�^�4L+_%(�|)�>i��5u��e�%?v\\	��7�P�������*�]�H`�PO!*�k;�3#(N���y�o������e��^ۋV�kf'�!e��ׅR�z�β�o���8[�"u�-Y6Xֻ@U�V�d-( �(	�&^7��Q�iU��=�^��q0�6`���&%O���Eף��`�Ӌ0�1����M���0�O���p�б�����{l��S#,�:�*��=J)por"�ؑF	��$.��2�H�A���E�<�@�h�0�t�������+���������?_�Y�n���~��Z�[T�b�?��C�f����^�R�Ʌ��V��賛ۅ�j�a�8��)룫7�Ϳ�={5���*��v"��#�"{a�ﶣ�FN��(˓�#/5��[��Mܞ��L���$0B{^^c�`�	���$��,#Q::�M]��I��&��8hoѽ|�^%�֧��_n|�@�(�Mlb/��|����n�J�G���%5bՐ���
��Z�T`�Y����Ͽ/�0��X{��״A��F���a��.���s�!ݍ{8���d���ǧ>0�G���J2�z*]�4>w\�]ӂט�[yX�r�G~�x�jgN�3\ȍq�>`,01;�凫⿙d�.j�;�>y����L�^Ϸ����ۊRO�MxVm�$�Ȯ'��{��$}�/.$��94��1���#�LP!������y_��C�2wa 4���Ic RrX�t� ����eR�Nwˤ�ߵ��"�/VzacĞ��9��Ez:|gw���Ge`TCg �&#���<�,��� xv���̌�2l9t�ĺ"��Gl{z�E�'�3���c ���T��ck�(�a�Իs��1ЦT#eYYɭ������fG�wv?IyH����/���lm&v�ռ�'�����R�*���7S���ϸPw0[����G��<o��A������>"A�b�Q��4"�)�"@a`�z0ۏ?�L�"��2�ג�-A9�|6W���
�hfK8fU��"[5����\ֽ��f���� �A�_��S�M�i�h/'�c9���B� �L�:�u=���ʞ�N���x,�a�=2M��*X�ۍ*y@2
/<�S�إ<�ע"��=E����^0���\��FX�GHP6ڟ���(��@��Ԙ��x��A�w�~�QoL����qm����e�i�%�MO�TR8?�D��$�����O����I�׶�	�b?x�(;�G�+��M�;� ������-�|A��	_���D�Y�Ri�aW7��U[;4������u}1p�i��CY���r~��mw��$���1Y���;eC���M�������G�|S"���١-Ri>t��y���F&<�8���j2��	��]:��(��iKK�@&�+�Ԙ��2;ͦ��1�nHP�.���GRm�j�}`��:;�aX�ᧉ�i�������7�Y|����d�\���/��9��y�ӦE�e��Z���r�n�*Q%���P��^�RQE��ڼV�_�_�%8���6�"BK[��p��&�� +�KբX&Yk���38�׃��&��Z]2�c�5�	q*�z��oJ�����BP-H9�>�+?ݲ^G>��螖���Bf�{����;mv���|��Q���IQ�`Lܐ|N��
��7<������Q^�`����_H�<�ir�$����&�u�󺩍"/ftV�w�B��R�*R�;�%����L�� ��v��6��6������.q�۪f��(=-;/�m�L�x��J�Ֆ��y����H���ǃս+�Ѩ3J��%�z���c�A't��ꖸ�@���g�}���n���?n�:�����4P�'��$�O�%AX�oo7(?��'!��%��p��8��S��ǎc���j�D>���dgZ 	z��j�5�'*�CX�Q�k�r�=On����` ��J\B�2G֟[�������-�&�R�;�bi�p�O%W�}����nc����ce�X�.��LQ̎���3�ժ�[x�i������^@L��G�.h���<�(�8b��K#\W#�h��'ի"Fʱ��R�S�~Tg���̉442G.��^t�\u-Q�J����^�8]eԗ���K<l�IPg�~u߯ĭ���{�G����^�f�(��	���{#�6�9t�2�=Sh��n�M4i����x^p�eQT��������+���P�7y�j���$���Ek����c�G�H-b�ܿo3�a�P��L+wX��9��_yh��t
8��D�8~Hc��!O��� �v��'�]'�r������vY7�Vr���ܕ)���Y�;�$�W�dߝzh�O	i�!\<��]�
�+��(��ms�!9A'�r��C��=?q�X��4$_#�!��q`Fl�]E9 u]_P	g�X��_S��J�;#���Ң�܎��7ZV��#��{��F%X�4QSX7�y��@q����\ʶ>��Ւ�r�XW���=�G�*�Hjj�zg�vyZ����a�
���4���M�]CO���M�%+뻎�)q�G9OY5�!�Jy�}~�!���� y�m��� �6Ce�$�9�sc��(�J�i)�w++4�+�j�m�Q~{��U7�zTk��Y��P�D ���]�k�1�@˷4KLoϲ3�ĥ29��K����d՞�NI�m��:��S���iF:��i	���j4���*_�֯�� �O�;N�jD׾�"�$�� ����o��$YN���-��'������7������������1:.�.�3)�:ZK�Q
6����U�_��V@��(+Xe���!��z�O�b~��p�6N���M8�<d����O���7����0,Q���y\�R A\�6�"����SW#�j�P��N�o���1] ؍{�m��\?��=KpGܮXC��ā{��d{Ý�^��J:����e�uL��烩��j<.����L������e=J��<��X�A\�N#��osʊ�(�7$�����a�w�9q]�0'���ݸ��E�a�bt��t��c����]�ƕ��(ϵy|�c	8���8�*==+M}-�,��Ȥ��B�Un��v�����)�PH8�@of#7Jn�I�T� ��r�pWiS�����J�j2�T4�V�()x�ċ%�7_L���	�Ut~�����"������s'��H�}����Z�։��˦����?���
ج��B�R���Fws,�eov�k����ר��:zv�^Z b:ɚ�kz���_Y���{r�d�<���B��l�8���DE7U�]�]��,Ȧ��)�WƆ�dWX�u�Oڃ��?��g����N� $ ~��������{�hP��[*���sq�}߮��N��x�;���4�K� B�Vt���d�#��/���*�rJC:~lQ?��{z>��*���9#��
�\���?!D�bL�y��6`v$lSOY$�J �(Z�@(�X�Ĩ���/����[,�q��{+
��DȔJqߧ{�
��K�?��0O&*u����&򧫌H`_JNʨ�8CL<^I�?�"cP��E��R,j�k<ȉlX�R�������O�l-�j�?VM^KڮW����иI���-���S
� $Mϕp����b�cJ'�����#�����7�E��k�U~��~�ŰU�q���X�N�d�7pkH㎌�������4�Ҟ��yŐ��\�{���x�.jc%)>�~9BwvEtO����jm����E�%~\��)J����鳚����w2� ����ȑ��ܬ|��G~����C��Ĝd� ��(ߖC,b����y�J)���~����z5J�GҴr��'��Ey��.��$����p����m?K�w��J�� �p�@��#���O4����V�J��i�K�X��qJĺh[�t�	������yXф-��n\m��y�?����t#F��B\bG��^�%ڇd�@� id)S��H7�
`��Ƥ�����ys�M��eq�6E�ph�k$�6��J2�����u)#X�F_��9�����̖혥�c���o�<�9�?T6���4[7\��AO�d�OD��vk�5��ԫQ-�����׺�<c���$��[N��9��Z���&I��������h�y��f���r7�F��z`7��.t�j�4N��O�l�����(L�n�;^8��z(k�y��2=�D<�"�����(������� r����;2X��_���˻Pxi����o(��F*T�g�J+]Ȁ��l��g�t՘-I��*b����@|u�|7R�]�[$hH��:����!4[�4������5Q��o���@p�j��R���h��v|�v0���C8����{�IVb�l�͕���|}�ٍͮ����f���i���XO�Q�#,x��D�,I_��㣵�Y./�[JH��3X�n0�VF.f��7$6�nV8h-��vŻ�{����KBAB�D��E�Q$:!z/ѣ�6%D�;�(�{��d���3�0�1<#'�s��~����g�g���GȞ����O�{����.�'����*�V�7
'��np���w���t�}/��:���� 	�ݓ�� Ң�'��ٻ>�8��f)p��x��Fdk��)�lTh��,qZ�"Y��_)y?���)�9d���-X˄���Uj+sYg�����z�F��f�@@��n��j��6��:�2+���Cj����(kf�`�:=�c��z���b
܃�K#'w�|�a
1<��jԙ䩚�_f��El��*�\0R�l��>�L��E�ْ��o+�&�mڸ-�v$	�ȣ��}�pV��ĝ���r�v��=��w�w�1��­|MՍܒ��6*�L���*�,A��#M�[�V<�) �����=�hpy�?�8�` q��|8�̄9�xn�{Q��MYsC��y��ɞ,�-Rͥ�>6�U9�kq�;�&�����O�V�,O�:������$[-~�@r��ұ���|�4�������/�1��g�����7��ꭃ�ށ&��� �-�h��9K::�Y'+�{�Y�.#��Τ�<{GD���W�5���e���7�%��E��p�UZ�X��+W�*�q3ۭ�٨�[5w*޶��!�a��|�{1��x�.�f�Z0�G�cRBc�]�CEr��=���|������/��qG�r/{o֋���=�8�M�g�v#UWs+j�&P�N��Y8���MɚG�֞c}�Q:ߎ%n���eP�ec����}�$f�g�P��b�r@IT����x|�2�'.d�S\��f��^�ɝ���AUՂL�4��7(�n�{䤾u��4���	�}S(]�!��E�缟��F��*8:e�x �AL�b,Xx8!m�y�P�=�lW����f�7}+(p�↭�\���=����v����l*�p�As��Y�*�22-�Yώ?4Gel�ɵ�h� _m�ß����r�=���}�ך~aGһ���`s2+%�a�#>� /&!��m����v触/��t�`�T%��w���s?��F��,�t��	>�-�,�<��GE3 3'��c\�-q�٣��p�/�Qv "W��C^4�h$�d�Ě��0��*-����O�A��>���K�����K��"[!��:����E�O�p�<�<��5��p�"q�mK����܃����3��Sς�Tܒ1�Jq9���N����S��-�{FL��Ǟ����e���ב�8�c�h��K2�|�@��^����b�����L���a����-�>����Nh�B�<^P ��f�B��l��gü�C����D�?s	OO�u�Pc�6ƺ�H%xZɑc�2F2�{',p��`2H"��jټ�F�[��
�E?���;�|�Ň���G�����w�k�g�B��6Br3n�6�y�^ϙ��O���ԗ�̙;c�F���Rc�����\ڨˁ�j?�7FA�4�?�`&iR����Z})��]�����2�WOu� DU �9i��k�WV�1��4��I�0-;q^Ϙ����{ax���6�kJ`).Ԁ��l�p��*��(����#�����ڍ2g.��gftIhLɈi�aT�w��3ˉ�GQN�ɕ@��o������S*0JF�۲j��K�O�W�L�T���K�����>�!ۍKT_'��f�M�]��m���f�\�����k!���غT��o�&�$Ol��u��S(%I>��e�1�k{��#�����,>�j���mL���
�-H�`��RLp�։E���ʱ�9%걯&�V
5D��=��A��-��Y鶒u�>p�mņ�|��M���;ɛ�SW�7��iN�ֱ�v��
T�����ȟE\�/f��!D�]t�)E��!&����YL�����Rj�do��k҈ǹJXS�Z=n"v��
y�Z�h�`���4��J��e7�G�t�G�#�i��S�����^��R�m(U��^�q��J^��.�8�=+ՄI��Œq�� �k幊v.��f��\)���s�Dӥ�U�q�ڤo�g���>�N�{l�oy� Z:�#w]�*M;�i�FS�0"�9�����-s�F�ίr�m9��w}b/�v
T�W��N7ip��`�:�A��]���JHZr���P�а���*X2knTi>�ֺxv
��s~R��d�c��tN�o��UJ
�e�B5�
:��%�s�V��4�B�m������#AX�E�Q!ʾ<g��`[���Po@*�*�����F��8O$-:�ō�+���(&��dP�����m3��U��z���7�ܑ}�A唙~��;�`���sf6����o*n�R��)�����[^��hf��M�蔯��o����%�Q%��X�2B+��,�ct{�O��xèKC5'E$q�vK���>�)�r����Dp������W�ҺЗ��>��wZ��5]��c�M��yɪ�#I�8S߆���B�s9	.�����[K��E�R��B��S;�}<4瘄w�:�X3V)0�xt���~�]���I�U}�Vp�q�-�eE��j&�#����k�$w��qK�X�:������{6��nt��/�1�z�E�+�u����P���j8���ˁ}Z��uK��ڴ�hEo�ߔ��fQϡ��K�+p�"��,y�nnm�y����B{��J7�i�)�@i<�*w�$��!2c�tÛ�Z�̉�t��>SG��U�H��wVڰeѺX�a�N±L�R@`=,Y�ýq�_p��V�*1��yJ���$�L�@P,�E�l��Wik�d##�!ϳ�%_��w�4����͕s\٧5u<ʗ_�C����u��j�m����͎��P��߂��g�U����f���)�q��b�א�ϕ�}���f���L�3m&S�o��*W��N.�z��S0�R�f��Q6��Z��$�O�re���e�ݡ�~�5�JqPo�ˑ�.�X��oԵRE��xp��@��3���\�+K�]�E7�`D���0eܲW�͎x�kA_�@����l�ͅ�۶-'8����(���6� �d�[^�c�>x�i���m��=�OwITq�*���ζ�㿌��H<\��Sl�%�3}�r��p�-��3����FwW�R?S"����RA�UC^����ۇy�=I��o��`�E�dh�?�n�[�iF�hY\YZqIK����[��s������5\�wז�q�0�͌uP[
�:���QB��E���!��9��.w(�
b2�'��/`�$�-��4yW��?�@���B�*���w?�?w����)��8h�M�V�Ҧ����c����w|�$�QǞmR��/e[|�v�<?Ϧd���<�Sߣ=�A���wKY K@D��LqN�v��]܃N9�T��R����F�?��_A^�͋O)9)�'�勛�xxAw!��x�2����4��+UJ��VK���tl U�0��uk��k��6"Pk��)i
��0
��a7�)]�q�@�s�9K :�`�OA���M*y�5��2�wA9���E��s��-�H{�H8��w9�Yk��-�������T�F��']�終qw~j'�)H4c���q���0;�X�1������(p��C�P�~�mT��n���*cwc8�G[�C3�c�'�@[Q��ņ�Э��c�_�m��k�^�Zq	�h.j�<�3�O�f�-.I��?���-F;�b-�%�O`�A�������V_^�nz2����V�wq
��k�_�Q�g��J�8��L��b����S:�I�%�AY>'�1`�)_\��r<�M]��e�����6�p#��+l�;96�V�:E�WZ�R����@¸�⪨���6��ŕ��Ÿ�Q9��� �ވ�ȿ^"�|&fY@�⊬"٨فF�*;-5�n��3i*�4�FU�R7�0(G�"�-N!�l�N�?J�kc?����@ۧ��_X�}x�M]�m�d��!�Y��SW���Ӑ��nن߱��<�Nߗh�`I<�8Tv$s�4�_3�\����?Y�d�4bw��"Jա e_\M?�n2>��p����_R$�^w iɥEݫ���F�<�-��C	�i��EQ4�Eof�{-7�	����=@Q^�h�y��oL�=�&y��|p�����I��u(t�(z4cz�ЙKv%��m�
[?F��B�I��ؘK,`1�3��.����#[(��#��j1J�;,1���GwY!�@(��v�3�H�z-��E�����׮�$�I�8%g���s�/�k{�B�C��[��9�>����h�~�ͧsψ݉ڊ�G\A$x|�AҤ?����v�b�g,�U�=���N�[�zˉ���ӂؑ�m���P��8� =6,��^8?�j?br�?�1�<�|�n �08�4�ѩ��2��"'P�*yT�w�Vnp�%��>n9�s�Wtu�"&�4�&�y��)�����^s,�WCe(:��#~�X��Z<�� �I% \ތj�	�]~��CRr�8ǯ����(]x��w���F'�ի��K;VƊ8]U��:쟭�n06wI��,Sq/
��1�Xq�D����	Ο.+�V��2��m���'�OJ>&�$���K�*����&Uŵ<�LШeY��QĬ�s86��H��C\�S�L��m��خ�ᜩ�1o;��܁�i[�M� 
������4A���6n�����V���2�T,b��B_�9ܼ�W %2�w�T���w����T;[�ά�C9�=���!���nm&t?��{���C;?G� �W����?^��@Ӈ?KH3��ۚ�%¼�����L�Y�.OzFh���گ��w�]4�q�<�F��}s�\��	��MX�����{����&Z�Cu-c�f���м�T�A����8��X/�8Tl������o:i���KE��oQ�^��

]0*�n7��t#u@e�@�5��4��z qt�y}d�Fp�� _���D@�
Ԣ��p�ڡ���h�V�\�O���|���-��`�d'�Dڎ�M�Ʋ7Ԏ���5����u�����d=e��?|g��;]�_��$֨��jol�{%J�J�b�O&������۸onTC��%G�1n~��p�Н��W_��������V���\Q�8��wش�w��۔��lNj�7j�7����p�*��%��e���F���n*f�5Ľ�T����nQD~�Cpu]�$�FǠ&"�������=�>�)ڋ/GX�xҘ�R�Ts�������Ȕ5�]���?4:	&ǫ2�|^Ѽ��#Pr���d����6��X�igמ~�▪�)����+��kf�o���u�g�_���8%�\0W^0�<|�������Unn�E�pD�{_�u��bU3�T�sVx$��j�X+����F/.�!Ƀ]���c�ފ]��R%dcF����t�W�7RR�R3A��j/_�����'�ԩ�)9�
Pqkx�A�v�^��ÿ��o�+N���2��?^:�~����ȍ:�� 3t����PךK�/�nȩ X���<�}�4op�,āk��[�O8���'?uv�zSޖi�u^X]��_�.?IЉ�m�^)���ے��ԍ�+x�Ť��-:����QP���p&俾||�S%���C{�FV�(���~���_�@r�/���4�Ő�ő~�,q�Ӌ�\1���-�xxnx�­�����/{���V%ɿ{�{p�@�{D���_a~��iH�kC�_�堮$��!g0���=R�`�{w�F#��\�/Ay_L��w�������.Ns�]���
�o��O��i���!��.M��6�4�V����P�QkG���0��?r�HI֪�:��ك��lY��R����%��0��ݛ8��8�ǹ�ŋ����[�����l �����
o�ߠ�>��L�q��#�@cB>|���,��=yݞ��.å��@����H�r
�ܴ���pz0=��j",�)�����7����۸���⣘�|� ��oZ��w�?/��Կ������y3f��֭���A�:��^���տB�+4/ ���M��ܐL�P5t���seBymd���_����8r�?���C�&|z$ߪ�Y%4I\).� �SV�*Y�|��ikѭ���wM=S�FE�6��XѮ�H,���]R��w�o��?�z�	��ёW~�-F��e�)�������]��I t���K��Շo�/z�u�_&��FPL�^�G��ڹ����zf�eyF��O}�OT��g(=�v�������8�c�e��D���ΑE7tό�G,Pjz>���*1$}��uk_�0���y���i�z�k*��[��3<�ி#����5!K�I�t�t@9�6xi�N$�m���\�k%[�Ћ����d��a��'ɺ� ���a�)2�ʒӉ��R���\&�F"�k�O�ה���EU���Q�?��7E�Y�O�'&����)Ț���&��Y%cM-�j����k�De[�	���Tcv���UJPv�7��i@�R�'^ϐ5��˸��\�,�Oh&��	oh�5gD�D ��P�y6	�����d]��Ϯ����f��� �\��j�e�~���K�֢�c����"�Z���P�Գ}*H�|sչS�M�}g�w��Rk1��jFl���yt��&��y��J��k��Mw'�ݓf����\|���{�%�X?u%c�X�Y�ע�B�;�4r��WI����n�s�@u�$�_�G�2��j�֭ěf�T1JV�*�1@���0sړO�K�\%�����_���2L�ȡ�+i����6��63��)/�G��Z'$Gt��t�J����lC�w�/e����	��"��>�3���$V��/: �8��حN\�Be"�?��2�{�[G�9y��g4\�L
v�V�wd���뮞J�(ň-�?T��s�*1H�NaG��[� ӕ��������g���7�y�w
\�e#���g�{JyԞ;���e�_�E[���2��s�,@ ���a�z�[.���l��{�r\��]2b7��������OYJPc@$w���|��:�Ɖ�i���KC>?��<8y���ݿ�?f���5��mJ{wz�$ҒXK��-q�a��O� K�9�!�*����B5�����/���S�n�����`����돜�)�[bI�2��Ů�ova�]�3�{m���܌v�����K8����[�d��h����+u�z�Ƕ@��ې��2�>������E��^�Ġ�"9Y:x���U�����Z�ޒY[��9�������^x��t����H��k
�S3����ߖ�O�4C[GU��W0��n�_~{ll�)&�ٮ|���,XM`�7�n�S��즡���L��k��I�3S��������.�aE����MB���ƃ�MZUCs�<�&{u���j�|n�谘���'�q6��H�?^�zedF�[����.R��dY9���'��z_�����o.9d��2��dh�p5�d7I>�0�|ig�U�HW�h>���Kp�L���?�`���/�F�������G�^����0r�Vr$��j�]o�I�M���%�tl�B���ٝ��ۢn�9=�?I�Iڪ��o�8SS� �L"C��<A������:D�������uѡ���t.�42�k���4���'y�O�Ths\�o����wi ��ի�m��.^<eM�8�{$&Ӷi�H7�VTJ:��f��#�ܳ-6Y?�=o����37�{^à���gs3�p�l�Uk�4�n��n�]N/�84t������2ZMۓ���Nm--���Z:!:Flp�t�x�L�	fg�A�e�%��N2�B8�x�O��Y��i�Zܗ(��u�4坉��t
t������]���4T���w&�7��7M�VM��c ���ٺ�S�nY���kE���O?�+}����$�c��t�;Q��U>y1Z� �̻s&H�@�L�G*�k��akW{��lnbK���I�%��&g�]��u�й����m�}�<�m@���}�{�y1���/	����[�l�Omo���t.��䧈���[��2�Q���d8҈˽����~mT���(+��z�޸� ݟ٘�匦*�d��}�;��D�K�������R�N���5�Έ~��m��1kr%;�#J�i�3��|�֩��I��̼�A�K��R� ��
 ]����T@��b%�?�Se�5M`��G�'f��vo	��f�_z(�..%�����a�c����S�
^�����R��|�(K�)�c��b�zo���N*B09�=!�7��<߅�恙s���|�g���C�P��r���a�7�NQ���m�OI�]h�;�i<�n�0^K��L�SZ��W#��Fŝw̝C��r0��9�F��E`g襸�����j2�[� }�w�ؖ"�7�s�w,�Y�Dl*����"�o}&�ܥq�%����S�?p庽��qq6�^���]�9'��[�=D}28��ϛ�	ϿJ�^�g�ʵ*�S�c; ����G4��5K`����(�麓ue�W�ӻj��ft_K˚��TM�t����N�/��"$Rwj7��@���\+~�XFR�DPbN�&LdQp��#��|�s>k�;���:n7G퉜����f<pt�^�{'�OI+\ck��P�ݙ؉s2��S��L�C<eON�٥:���\Jk�z�x�+��i�H����c��Ƿ�3����R��T�f���l5p\�?9.M���v~7�rS~*r_|�UG��e*���ꂉu�P��������H/�`��Q�ͩVY��ƥ�v��G��dA��F���,�{���>,e"�3h���X@��y�p����}b��sڡ���IOS��JV�d��Zm�?�^�{ˊ�y�����[�������~�l筫�W=E[�Ug┫��A[7��*�'=��.�T�X;��]�S����J;���A��"H�he���	N"�����yM��޻n{���e���;�f�[Ug�
�q�=��q����ڝ� ��Ά���s&ץhqW�n��YK"FV3�3H�^�*��8�_�0;cr����Nʿ>���4�H��K��`�Y��KD�6�Jթxs0�B)~ޠ�AB Z�������'i�,�O��|�[i�m�޵�؏�&sB� r3qF�Y|Z h滙H�c�e�,{�������s;�ɻ��v�����s���L�H�@7����. @z�X7�,�����z�*W!6�O;�n�Ԯ��8�Ӻ�!�ш(�S��h��qT-<����?�R,���w~s~��!S�.���U}�K���fLǫT�XU�8��{Yk�"7�F�rw�_��H%��gE�>y�E�i���Rz#��K��[����TR_���F{�	-"b����?�N����QU�R3���D�׏I:��Vd�,'�Z�XY�y=a�,�>�2n�?��]�.��iv%&��I�.�&��`�R�m����Bn�~�k��I��LG?�|�	�qd��C*`��nd��+�7�dz~����UX%؉"�ݧ����KMU��w��ț�pMc2`�l4ǭ��0ʩvA��ϡ�ݴY�1�dbV�~�#��\P�/��*����E�
��ܲ�dn���-N_8�����eFX�9�d�Pb��m��%��ր^�p��f����>��"q��DԮb�"���@#:'9��A�s%7�����9ޜk�=N4�//����$���+?�#A~�b���t���2� 	����(~u����@���3���U�/���y���+��hL;�C܏�m�5�F��A��%�1uo�0lE��׻�3��!z'G��L��d�ނ'�XnL݅��َ:1�:��1����Ƃ�3%� v痙�%���yo���b���������M��	�|�y����\�H�=L���'إr��U���1R��e��� �T��7Q�Q��f� s~��բz�g���ҏ_�ᬁuؑ��qRb[%�\�����K\pZ���$X΍����""Z�x�ַ붙d��p��v�_)x�	v�Y���|�y�u�����-To��L.���}l��lL��)�&����aA[�H�i��Q�viǶ`� ��R�A���|�.@ܴ�M{�i�5�d�dU�������mt�����u+�2v|L�6��Nlnf'`��b跥5|�Λ�v�n0d�}`#�05<�~�D�9�i��ì!9�u�,*64�*L�l/h�p&�ϑ�@$��g�1�m�&Żm�������^l����m�����`�4�cC�#\;W�UC�������18��@�-�*��m�:�vp �ON���N��������K=����%!�3�_*(�[��D�V����"�(�m(#�:��./�ER�s�{�4��K�����FG��5
�N���Y�{�^<������}��q���0z�d�=�[h!Gc��ЎeA��i�������G��q�
8�Jf��$�������	����)�B�b��=X�^R��a�	6�(���&�vm����Z����2�����6��V� v�'�u%/goo
�ݘ�ߝ�PU�;�^5�G���w��[ї�!�ka_
7c�O�St�)�g�	�1�^��c�$횁���������k�+�&aa�tG���X ]aL���e�����c=өr�ݼ�n�w���zP��횵Dʨ�/�QR3)38Q*�	\�}U���(!�b��L.�sFNH�<�/����*�
)����d�����.(^���Q�ܮ�[<d���gؚ ̉���n�с
2�PM��{X���0]e��Ӡ;��ʥ�� V�:m�iH��h�L���Z#�S4}�Xjj�&�Vۼ*Eu]��#�u���n5^�0}�E�V=/"m�{xh����oKmxx;�?6|�,8D@v,��N�v���n��?�͗����UE@.>&�Y��-?>u6
U~-��l�� 3��Y��eK��_���N��{��yO���@�0���&�w|�*���֨ך�yWGQ�N�����u�n�n~�I�!����������,��Ð�[N;�����^zi��Kb�û�F�{c�+&h/�d\��Ű�����qx�\^�.�����e��Є$�ߊU��.do��҅�V��dP͜Ax}�R,]�VRQ*mt�ѕhE�Za���[�j�X���������_vvj�3�*�tf�ٻ�� 0��_z-�*\)�e��k�8Ͼ䄖h��g(W�0;\�2)�TϺ���ׂ�霰�)�ـ^�5c����`Z��pD)F��P+�z��[��5#�A|�M��{A��^⍥�('T�|3��S���[�t]��_��N�ݦ��H�c�=t�5�i�u�Qٚ,L�SV�~?k���^�!�.��~��6�_�ɗ����I9y\�X�/�r���B��f����.5�o����g|�c=�.��$T����q�m����I���$y_�����2�����b=ݺ=X0/�6�Z��+��2N�bN,m�܅B�wS�V��Ɠ�o�w�<�a�JF��r�Z)ǆ��{�gc�3OH��? ��;wTq-��D������%�8&{�	�c�p�h㐿<���?�tqY�|hn�+��ԕ��HhF��m��j8�^�IR(����s�ĺ L:�[�c���ݜ�3JNىfb��NЂ��ٱ9z��]|�L@�h�z�u�WP����J�o��H������eN2���5��:��*-v�e[��W��7�ϸ�ҳ��Eo���E��H���.���A.o���O�C�s��E�}�h�M�_L(���Nu�"�&�5֟?훮���}Z<�#x�q�d~*3+f� � �,?c`�Ȇ���(R��C�xo>#j�zs��>Nݘ�U5+w�Ml�t��-�Հ��N8AK�jp8{��0�R�c�/o�+���e@Б��
�tŢ�ُZk�O������
�n��9Iާ\~*�yw��7�L�h��_c�{��W�Mc!kreg�|��`��g�
��΃8_�o����Y~�7md��v��x2����{\L:�g#�_�u��8���=���`���u|P���a[��ʬ�Ge����s�%�>�0!Xs��������D�IOT[F*�o�0(����%wc9�k�(��>����}|�y]�+!�_9�b$��od���Y���G{@�g����4�xO�Զ�`j����1c?ě|M܂�O� <��SbM���ΧU�_+mF��|_�i���	{����Z&���<'VR��C��=�z{�!�+��.���)a{ݾ����i��U�sĝ#�pS�X���0�W���e��qb;�m��ʛe�_/�S��.>�/����֐CX%����z�[Zç�!�>G�~u�����ũ�M��餵\_}A��-H��'R��2w�x�i�}=p��0��m���@F��/����}6�~����F������n��9��XŞZ�ވ��kW�b"KO�eUlN"f�ě@� �q���ͭmvGYAX�xF�^�m#�bgW���ߊIG'�U�Z�����5I��Dz; ���1�U?۫F��=�_EE��6��J�����;��U«ׯ�o\{b��*�-pʴ)�3Q�K�m2�WP�'z�}��'��Z�ݮ��M���-���H/���K�I�zLF�yAy떾��5�v�Q�׼I*��� ���c?2�db�R����fwN&������'�9�{:���S�s�^wԛ{6r�B�p)���g����4v�6X��F�0&�S	������M4�|V�{�����($oę�@u�=Ǽ����8���z�|���3p<0}�����K��m��	�PöQ��|p��ii}=��g��[���@�ޢ�ީ�zթA/�r_�޺7�}9�1�T��v��7̎��ov�pÚ�S�P醾���Y�)�%��Q�s�g�#HZ��d��o6,N^������.����|ek��jU�� [[&z�D��:�u	x�l+�+����鄗�|>��E$��e�H$�v��$�)����Um+,�/'�9�E�����+�}Et/G�����dԻ���7����2����RT>�?r��lM̅g�b�~�����}�I�_�z���G�9�Q��_�2V n�����(��U�4�nQ�
/��k
DXE&��s�X��N���Ac����w�"����2/���jJ�йD� Q��+�q��� \�n[���xw'b?;t=(��PL�fX4�n��k	q!��9�\��ߐ���|�Y��P��s�/��e�k�g�5\�|l�sf�0�k���4m00�] ��܃���rt�R��	��YQ����q����׉/��WR�ڝ�D�.��$Wب-Dl�����7�������H]{ZK�<������7�z?�ZDE��q�D�*wo�O:�����v���Zk��w�r�2�V�a=hLV���{e���>��@љ{��L��,o]W0�xR��i��gg�����VAro���")��a���K�5N�g�r��hg��r��k%J�IsJK�\'�M4�m����Y��֎"&u���@�zbR�i�|b��@e+�H��#��#OUy��&�N�!b�����F���䭛��lL��Bay���o[������d�����������Ks&6	�Ef�ܰ����A�&g�j�~"j*��>�"|9(u�)� �E.� @FRo�M"���28�)=y�0��	�*�3eC�9��yWϔ��k3���x�Y;O`�x��*�={X��nb�.b'<��jkd�R�!���q�������m���k�!J֫yށ�)�,�v2�*'���s��Lt�[AVVKmdR��!�����~xs23��yx��iK���WmPid��)�c.�%�}�$ǫ�����>o��j��v�ɕ#�V�
�q�
(JR�Tk��D�ü8�*+qC �S5K���;�����8a�8�*l��vz*��#L�PYD(	c����\�|�,R(_���x݅���d84���9�֩x$�H,KN8L/�R��6�;'ϭ�y:������<�S#�Z/B�����+6{=ھ�|)�u�^>�d�U��H��KrdK���o��!��#�p��7��ze�yh�"�'�������,V�D4/��W��Y7�z����t�t����V+d [�?6�0T)ݮ2�RYw6K̰_���W���,��|ˣ�%W�S#�Yņ���a�����p�w������ZK�j,� Y����*�u���<���t�F^x:o�w�d�ڧ��d�͑[v�K��x�`��Ln�~���"��r;��k[�;곱�r]SL�<n�ie�z�#鑬� �?�5��O���pQȮ�wC�J���������HM�B\�{��ΊY��tӊ�x�E=�#�G^r:1��x!D�[�g��$\�Z-]���J�φ����8�<�4��	�9*&Ψ�AҮ�Ic.0������)�p8�N`��U)�!{�E�Z�X�C��8�G�2<[�J��_���B��G�~����|5�U�ZoWm���Ҕ�O���i� ���O�^�c��i'?��\�v�q:`R���]� z��P�*�<�Ⱥ!ۈO��
H{D�C���sb�j�os�A��PwgY#*���\��l��Ul�ya�'y��{�c�F�_������x r퐫�Eu+���"|*]6���e�Z]�#��@-�}X�[���z���ɥ��#�!'i}�|�T���ɂ\����H?�E :I;��r�s��Bˤ��>$^�1h9hf;Q8]m��Xr����%**@^�ϋ���on�bk�Q�j>�)��h�@a�^��W�6���!��� >&6�Y.P�-U�i$e2>��.�NܿO�P�.,'���C��Q����4�5, ����5�{��!�{��oƿc/���K49�]���8f_�{��M�,���9��=�@������@���Ϫ���@��G��kӥ7H٧�_�,��.In�������a9y��AV��.�3�*�;.��Zݙ�c��<	�Sc�a?��Ո�t��d]I�MpZ4��E6�Ȁ�}r�d��l��Q�[f�Oͽy3X�Vldf�ɵ�
w߿�����6�Kzk �WE�~�S�Ѝ_���\��������mg^����PR��!���3e�۟VM����D�5)_�E���6������l��@���7ԧ8J�G��Q��9O��en�ܯ<�?�/r�Y&�Xlv&�Вs�W�ה��a!aur���k堖T�@v�$�#��]�!�x��O�Op�m[���5��0�U\�̾�˪�7K��u���S��~�{[U[�h���SR2b�]�bo�T��cx��!�)d��������Zbzf�}��sw䱍��(7�֯%�����Z�9�$X�����"�k?��W����� 篋���χ�2���DEG`F�R_)���y���y	Y�À�vP��'oɶ2���ƀx�Z�˦�K6�!_��Q�e�|���ޚ��n���V̑�_�G�yvr~&0��@шظۀT%G�o߄l�6W�{��=�=�>e��))�G�~��.��4�3���3 #�WD"G�Ѿ�����&f|cƠ�/�F���U���ط�S�����2C_*R]�{u��o���9m�1ȩ���io�y*�� J�Ye@�6�E(��iHS��8y �^K��N���*�Q���fS'%����H�x��[vx�ª�TQcLíӦ�u�aC-��풇�b��=�+��"�ck�s� �5��L�M���[���3\g2����{H#��VBt�Rw|U6��t�,A�JJx>���2�"~��T�R_������^5��eXY1���<Pt��%���O����!��������{G7��0��O���)N�������S7r�y.�E9S�}b8��Z�,�h�y}�u��^k~M�`�6�����D��bt��9����R}�Kzy�wב�Q�0�A��7�&E���Zƀ�$3輸�~"ցJ/�n�F/��A�EL	��H3h9Z�Fp��*��3sw�_'�5�?�x���c	ڣb�9��c?��JX�]��TRup)67�����yiyʦ��z�b�醶�����ܭ�|��k��kq�j��X���,�G�g�Fj��>�ICj��&?Y�R;��sH[}���ƙ��T9}'����1y��hת��U7u��$����I_N)$�.���1N��BN:{묂l����S_-X� ������r纖hB.���
��,�V+׫��F��.�%��\�V5�t7oF��<�(�9����x����E��B�/����rj��E�����!<J6
���|��	n�IAq�m |�S�_ y)7#P~�ۏ���;~������&���b褽�
�x}v;���,gA�=%l�Ŀ�LÐ=�`kD�R��+xM�+�� �k44x�
�ɥ"Z�[���r�<+n�Y���[�.����e����-���@ ��o�1z�ھl!G�y�0� ���&����/1��f\�IH�M@��]�G��ԏMx$�\i�nSM��Pn�iv�N�녎�c�%?e~Ҫ�*N��&���W�*z�#������z��Z��Z�����*�Eyr3�9��Q'�$,9u���}���MmG��]��=4���%�E�Ʈ�􄾹��n;[������]i����,v8嫉�yHa:pj�M����K'��E���U�s��:s�{�YK���֭�ukF�S ���94e���}^�}�1S��SA*VN�sT�о�QlH��ܡ�!�[����!�H�<�o�Q��U��C.v1
r��~S9k^�<�U�QB�-��D�b_!�O.�P��r��vBm���)?����щH�F��j���km�tY�R���� ���ڇGPR	AR���T@����S��niJr��;�c��a`����+�������[k���מ5���teW�^fණ�I)�
�柌�)ƺ�z��&�|kň�h���M���@�TXQv+>���^l�����m|u��"��ۖ�Ďϖ[�j}�fӳ���2o�>+�������|�&"����͸��'ݩ�3��ΑbQmפ��KD��������0ðׯU���r�(s 0� K�q�6##������*�����$#�OIM�JN=�C��GחOV��hW���HZ)QP>&/����`�tHZ�[@�_Q��Nr$�dDl(IH����%�-�K� %8�C�[�J��U2��6�V6��_{4U��%��Bkd: ���2��j��w~�lƵr���|z��)����l�2`K�O��3iSp�ސ�Ԟq̈��.��p���(�ϼ�k(�-P�Y=�k	��+g��+��]���	��)3]���쎑K�|J��y\nh���c�₭9\�o�)jD�ՙ�Udl�O��;I�E�~|;f����Z5�9K��oǋ���'`?)����S@�O����@�S8�~v�D}�J�k�Srrqww�^%$}�P	��o�I���z�[�*<�x��/}�S�j
~S��>�Gd�fٞ�l�hv՜���G�*9�יmGK� )ģ�%[�O�JFy	H���|%���c~�X��yˣ/�>m��|�X�!5��Yd�%��깿��rVt�u4J9b�w]��NZ��p�,�s 4�PI���쏢�*�m�����?�1"��|&eg緆M%m'��
+�cs����������=��'�w�r�x�&�i���)#C�s��|W8��v<}����d�DO��@7:��Q���Z�1�g	d�܋1�J'Cx�p�?��ѱ%}�v �� ����U���,\;�-�l.n���Zv ?`�"��ܽ&�:�d��3�Y���-H,�q�?=ԍ����J$���X�w��y�����p��kM��{���\�� ���0=}L:��`>Z��X^rvL�4�-z_ȁ����p�íqdrz�Y��.N�CL��.�**s�<{�፟_����F�x2���		�!Dr�v%�YT"a�p�����R���D.y���*G����ۇݦ]gK@�d����FU���l��>wV4��`s`o�����4�e�'[Y��ߣߔ'�z�C�?�u(0'�L=tpz8�v`�6�i:�'Ku��;ҮkmD7[Y0�O����M��2E�1����-��Չ<��/�f_L��&���e�j,�*�n:��er��9��7�
G�������rg��0��뎙�����픏�|e ����o�?��A��"��ɇ��5H.A��!`�I�d��t(5P#�2��SSk�&ѫ)L+v���ӄCr�w1]�d�.:?���In<⡦�M�����	k>���5�|�F�&�(C�5Yr�@Fr^pν-=��������c��?�g�<BN���o��-�?Ƌ��Qf���o|�m�����o�vFhp��|�R�؍\lX���������d�K�Q��m+��_1�$q҅<��ӘZ���-�1� ����p��o!<[](æ3�����a�ɟ�(m���ɗ���܄�E����}���c��vR�"�'�5�/���?����n� �&(�H3D�y#ʃ�WQ��Yɗ1�0����/����)6�:2e�	��.fY �N|y[�/�^�[5��gbN�V&0ok�6T�C$+�@�J�W�Eϯ�)����]���mN��~O.n��~S79��1����f�!��D@ ��p��>!��zY{��[�����&x�/'���V�k��Q�Td8\��b�Oxy��~H���f�t�9��n(�+�W`rF���@�!�b�P�)�^b{ �GaL�-��N��F��b�S��1�Z�v����3���699��5�RP&�p��;_#����o|�TM�7_��z��)����G(�m��ֽ&vR����^
�LLO�5�Ь<�S����n��Z��3jW���W�l���@��Ψ׮3w��J�k�?B��]H�枋�WG��4��Iݧ[����� �����Q�_�%cӌWj�����!�����u�v�%2����&��"��~.�2~H6�.9�aW'Z�~L'b�;Zr>GC�&�J�/�w~��L�;:�Hj��}<����9���K!:��¯���äA�n1�9@��������
�)���]�R�%���K0��g6^�����x=��*p4�]�2��i;��2"(;Yi*\�׆W��^V|̤��N��,�q,n��~�mH�8��H�p��r4�<�;�\�
��7m�Y���t�ɦ̰��E�S\w�~}\7���S�\Jݑ�o*�^Vu��.�v��M���O�:�P�������O����Ս�|��TE[\�L\�N8Ƞ��5�h���ì/��뜍��BE)�װ��1A-C,V�rѽpxa�h}bc�#j�q��"�*?etV��yV�D My�����(���6���O�d=�i���<��҇&%;������v�|~ɵ��A�ށ��츛\�U��,_�u�t�l�`�y��^���s{nA��ѳ��O$�����$���=e�}�,K��=�*���~f�`+�io�tk!"�?G� �D(��[	J��IDÁ��ٺ��]�g���ri�l�;���E�;s|ő�����Y�����2#d"a�`'���ec1���B���4�3�Ȁ�\��lc�b0�v�Z�2q������8�א_[�
73�#������c�J�-�!���'���u_!ӜUP�J�ڮ�8:(���\��B�1�g�zw1C�'J,��Y��+ѰM�-'�VH�Z����J���
x20�nh�B���]42�)�v�҃��h�ە@�� l�s�_.�}iv	&:D�h_�p�PT����)+�T�p��Y����?�F��Rd�6��R��cr��[��DpD�&G��I����-GZ���C��!�-�e�/o��D]81ߑ���� �+�W�Y�56g��`*cR�g&]]Sg��O��}F9JP¾|�U�[2���ƃ�c�KĹ�Ҋ�E}cezu�	�_��ɏ�]ޝ��7͛�l3�{,ש]�,J���ߦ�>�gXߠ��D�Զb���L���(���-�� ���Y����ڳ�Wj3i��������H�c�H���7�qnu3�|�ւ��/'kM7c�MX�:P�\Ø<}҄�X�P���<*"���$�'؇]h'��Z��H�>5��	,������i1�.T|=0�+7{��Ӱ=�$[zջ;��w�6S��|���%\�3bqz�'�r�(NY��Y崾��z�=Q`Z�O��pc�Q�ȯna�Z6�����U�D�4+�~f�A��2�E����?�G��!�F�f��������^V2�_?��8p'~�����W]Brv渚�CE����_�ۥ*��|[b�H��_�p���e�|��P^�����P��Y����0����*�� ĕ�hH�s=	�>��/�R�1���&Y�|N��[�;�	ed��p�̝+����y�J����|ӳ1�_. ��K:v-��b�*��o�aUKs��5���ry܆�Bo���/�m�M�,Y4�B���ՙ��q��퍑5X��&ЪL 7e���ֶڎ6k4L��]��D��K�L6޶��z-HEѹYM�#�'ڂfٶ�;�\��r�W�H�SQP��bb��$T�)�?L�n�I�Xu���9V5/����Ef��#0+P&�O����<�9���o�c���W��]#�l���潻 ����Y39̎P�4y(ʆ{������x%9�v�a�*0�j-�L�7�Զwxo��w0E$R��<�K�
s��������ax�xӖy,)!�����"L_�z#�ӭ֌_��ٰ������Q?}?yr��9�SC�\��yj�|�Iz�P8$�&l��F)|��"�//y���(�M4
~cjjl-Q2#<�$w�#��U�d�Uj�UA����� [
1e4�[���?ⱽ�~��l���8	��7�[��/i�8���AZ&BC̛��<��ꚝ|�+�
�Y��h�-u4|���O�PG�����?g}SD?J�"�{@6M����Ҫ�	����� ��ǁ\�ZY��c?؆�]/$�&�{����l�P�u��1p�Đ��kY'���]B��w3�(�%�;�7��X��̑u�1�N0w3Y��!j�.n�;���?%Ec牓�kk.��^����E���W�m�Ѹ��wo�曦� �����϶��5�	�5q,�2S�����s�/����|�����4��Rp�/V��2�y1u�@Q@�����pp�p�ޣ\��j0!�Ķ:\@.05Q�ނ�;-��~�ʉi�V��7{!�i?&����=�5ۂ%^1�=�V�8��jԃ@�k���Pm��	uRK�Bn���-��?�he]�(t�8s��Z8���d�:!Z\օ���H�}�`tt��f���(娊ʥ�J��|Է~Y�ᔞ4�'^�
�_zq[n�c��XX�~�||��"!��5�*{�VL�c-7c��5�^��;:��ڈ%�aK�s��I�e�%��S}AR�R1?��[Km9�r0B�p��U�D����	y�[����w���K�؁4bL�گ7�U�[���!��V���12K^��tUQ�4O��U*�T��fU�{́��A�c	��q	�o�ެ�E��U�LF�y�_H�>׃��s�P~Sxn�~l ���*�LN����ȅn��	�E�QMr-���o�W0�o[���\���VY2�~�B�<N�o"Q�`�U_H��OD-1��$﫩�r҄�*�!x�������dM;�Hi��M�o�Gl�yB�2����R���\M�������\����'Wxֆ��ɩw���+���m�����^!���_���<c�?�9Y_+�������S����My���~ŕWRzs�����  ���f�F���,������;
]����)=u�)�D��ǭa'b%�Bֈ�R�5���T���N=�L�=t p�Q5ð5׺���DOD��K���t@����3�A��Ԡ
B	���2h�ʟ�G� �>D�l{��.xR�+�����N����ßN'�Ǹ�E�R���A9�������yt�!�_qE���҉}��Yv9y��;��^\��n�S�� ���X*��r��d6���{g�����\z ���4!)i̳g��2�(�r:��)=���a��7j�����r�  �'�(ٵ���ۨs?����B7(�kd�(M�ma5l\��z���̕ �߅u���◠�z5�E��3�K�_(��rAGJA�os����!a%~<uvi�  �� 9 ���*w�O�ʦ���(�va���zZ+��%��E�nUޛTSb��.<�*��8W��fP����Q��a�miE[Ҹ��́p��ʇ��7�W� �P�
�L�����՜��$�Lֳ����$�q-�|�c����ع_/W2��;��#��@84���+6:[Ţ(U_]�u?����
�} ����^ں�EQ�N��PW$����UH��R�6�H�]?�M��m��K��[���r��8��Z�il�p�.P@��C��ɴ��;��@�p�"���(�) �T�Ȕ�$�R��Uo��"4�Z~�I�H0u�o$�Z�M7�� P���C�g.�s��S��X��0��S���]�)N�K�x�4?��[��6o9�q2�eV�Gv�ƩC��n�6j���ܵ�rQ�-�����$�F�I&�U"�f�+�,��N}��e��x�Jf9�5*
�8s������]?  ���e��at ,hby�-&Y��r>W��GW,�;�,�d�k$�޷��!v\e��S���q6~򇀱wX{��'�J}����~�*'��.vNޟ�,�3�RO��T̏�,=�o�� -�K'J��s��������(ըI\�����B:��<�zt�yb����T���@��:�Eh^B}^���sQ_��W�����/���xH/6M��@��O$x��F۔%��ָ��[�9cG���7_�!��|)\��\t�x�c�p���A�gZ����u:?�܆(͔!�wۃh�n�ʂ�s����*Hy�m'��ml|����noҷ���eJ ��n]`��z�[8�p�c�?	�XJ�#q����Ul7W�﯆��.�h�M7O�MTZZY)"R7j�=aL ��:L�p���}Њ���槼ը��	W�CBN:��!�xiB��1��&>��+��Ua���=�x��x �	M��4�� ���t:ޖ��d��Co�V��+^���ӛ�\\Q�I{Y�{�&���bB��6��#]�D���V��T �`l�(!�����R�\�� �1�1���v�E��%w��2]5f�B��u��e��^�>"�b4���h���[N����D)��� �.��'�I'@��0�����6/*5�$?����\���Y�#�H�-=����� NE��s�K�(�]� q;匦6q~�n2�&E�]~땕�ڛ�xD$-����7_β�x~���Y��Z��A��O�ɛ����,�s��-j��B��4��m��ԃ�aoS��J��۠����ܲ�l���%�Xز��w=t'ݯb}�(������}Wf��	}KY�+�>��h�>x��_����]�
}��SW"�]rC��.� Ȉ��'�v��
��ٴ/辟-	�����;��ԍ��U����c�q���+��0D��7�G�g�!�"y�]�g��3���M]"�b�7�C�農�j�ׂ0���{�f�>W
#茂�7��龫��8�Me�	_��wώp��R���9I_�4潉���p���@�T�m̜o>6���v�Y�h���*�W�\���!vd'��;,p�Z��+8�]��<
7���D�3��x�l��N��/s�4����[��5?@��U��z[��>��#{�"��x!�k���છ��c�[�j�9U�&���$W����%�@O�8&�c��W~� bF����n����ƪƆ����vm�5��lN�T ���ns��.]M�k����{��:;
�V�М��n���em3_�y�I���4kcn����2y��Z�$\�i]�# ��8���<�#o#p�*�2�a�ȇ2����\n�6W7�����u�쯓��e�'!�6�7���Zg�,e�?S�i��Y�z+z�
��Vm��?%S41�蒪����9:3����@D�����鐞n��s,�2.���N���UX��"���8��k�f�U���xf��c���|���T=f��㕌��b��7`�8v9��������GQl,O��4ld�s�Z3c�/�Hqg0j���1�e0��as�:���i�9�I�ϗ�~��å����˞(xϚx�J�F_/՝w��ߡ�I�F�s�﨟:1ܪ�� �=cU�-�z|b?%y��jm.�g̜��t��W�#al�����dE1��0�A�Q b��J���ugT��"O�����e��+_����n���q��po򶒝Z�Wm��X� Q�CbN~8I���nx^ϭ�Z���B?���ǫ����A,�[O�j��	E/e�P�y(���ǂ�S|�"ώa�)*�S>�Hѱ������MC�&+����,I�SO�2�̀������칑7��6�7G�R�cfJ���C����X�)vK�~����$�#�c:�G�q����}�	���Y�QI �g�b{��D�]R�]z`�\fK�!����'EI�C ���_*�b��H�Ao*Ф�S��آ��uB)���A��
 Hn��w��cU�y�-U�Z�L����h�ߊV(!�[�]��h���>U�0��y^�kzt����t=lWjtuA2���ξk����,#k5w��n�z�	���qD<	�/Bv��w�-5�Q?�u&o����N��j�]�[�M���"ӄ��-_c��[!�����m����J�<���?E��(�Ɲ�5	�hZ\��1��y(0>��g 4���l��w��  2�v��޺ӎ[BOm�2=�&����O��?�˻�C*�wf�QJ8�e���hI��Y݇ˆ�5��1��|S�&��5� S*r#����_{LcƮ&�Ve��֖Y�I��.l����4R�[�;��h4�j<Y?�m}�t��@WU����c"��eP�M����|��6��/��{GT�1�F�|n�3��5��[SGtB�;B�(�^�%X�	��_��,f�s��b"�>���V�X��6e�P�"��x
r,Q����P���~�J$�ɫR_$���@y.�e�(a�O�wU����$�ԋYwy�p�>yD'z�e"�V����F��יy�^WpO��J�Th�Y�T^n�����Vd�?s�������Z.�\��'�T�A2o�6�G���ה`��r5]'�t�k����[-��|�fMLA�����Ŝ�����o�K�����.Ρ�
�TOx�oF����C�bP]�W������u�p[��rn��S��GXi5��`�+�m�ӆ��6l�H�u���|�E�J�{�)�le�+\ꕩ�*o�z/���y�3�� ����PG�iEκZ����[�`�+h�!�}:1��o� DHL�"�ŉ4�P����
���do	����	�'^��YY��M��cu-��Oׅ�`�97�hJ����Y�E�.C�I?�7
P���Q�y����;���W7�!����8�B�*��n�H�	�G��Wy\����͓|㡐�gi��&���9�\�~v�ۍ�����f��L�BǷD��7�����z(��Ex��尐ʩ��tw��6J��As�'����b��j��6{DW��skE�۳��O6�'DO�E��I"]V)0v��j3*��%v8�߈�=Jn�T�'%�.ADO�1E@�~�v��S��	��{�,;�V����qPiey;�o�K��\�P�N��"p��5��>xq�o�w�2x)��~�׵4C�-�t���h|F7��	��ьI1�I��'��$a�ߵF�س~eA|帹�T؇O�f��mp�6��	�AE��;�����T[t� �PU��S'��7�l��r��m$�C=�LS+Q��=�Z8�7s��Ι��/>�{�O(X�&,�=j㽋�4o�M��|�o��*�#�]�䇳���;)���,FWUW$�ȺW�d�3U+���̫�v	��6���*r�Y�������eB�&���6M����$>H�ݺ1SC��,s��B��H�jR�kA�=e��}�d�qW�0;]����W�js5���"����y��؅��n�kZ��'���	W�v��
-��s0��E��q�D�.d͚c)x��'c�	�*�,d��%w��*�;�xK�U�76��u���c~T8��%|R�D䄇ԔB�<���d_��f��UHۓ�5�slC���=�	�0Mq�O�cT�'M�$�So黫L	]f�2e�����P!O?�5���o��*���߭`�\�g����Ye__;�H<6Gة�,Ļ���5o//j�k@�#�N�V0������U�X�s���~fbǛ>�u󏊙U|��9��bgȲ�qe��MZ�\!�Q�V饽�Nn_��M�ަ��̡龪�y-��1�.AO�&Lt��ܼ�CQ��0ڂTvr̀�o�r�/�Rj[�-��n�鐘{�5̂z��&�F�g{�4�:��ջ�c��`�N�-�!q6�UZ 
�W4��i���q"�,��P@�������W�_Zh�$��l�˕ᐳ�r�:�v�@z�ؒ�\������!�6΋hwl`N�iݣ��+⼰ȾU��y�,���`ui��vl~>m����Ku[X������R��[jQx��ӻH��J
ۚ6��l��,����KuD��'�EaM�!��|2�
�Wk�;����AŶO��K���8|��9 ���Ua/q�y�"rT� ׳�E��UZ��C�K���f\�ު�|Y6��h�N�@D���C��Hv�V�h�2�O{�
-1N�7��"��+@X�F\e���l ��y�B����
�1hC�{1��\,�
8��	�H�J5��vPw0��}�����x�}���C���C�b�ꅺ�v���
[ljv7K| �p���1qx��գKuCA-B�F���O���}{}*lZ��F��6���2$���+� ��n���!�+	�V3�EIxȌ��mi�6<H��]�]'�
�,�Ix&��י��N��8%rO���t����܅�d�L�4;Kq�.O<�t��V�����:,P�\H��;w��ȿ�cC�j�ww[$vMA����?�I��&//O�')�x���0 ���QA�m_6�>�o��Et�ײ|bN�i�l,���k�t[��X!��S�tG1�ٛ�안}�	�'�d��Ϯ�g�KrB�A�Ovvy�9c."�d=���1��;!ځL_GoƱ�������Rڋ���u�8?� h��i�|�:kS���>\80ڲ�6p���ڧ��}�]������բ/�/�S#xc�a�ox�8=I���)��ɷ��\w�7�8�P(��W��
��m�\��y(�8W�5Wu+�C���b�3�%��yk��Vm|bn`{s�t���E�9�[�@8Wa��OR�	S�	���)���m^[Sb*:����� lp^C�8���!�3�T� �3�	����n�e�,ݛn5B�� ?�� �zrP/K���h�4H�{�y�(�~ԅ���q�tY3M���|�����ݪ���Ma�/Lj�u�Z'!��lU�����⡽�%t�HocV���]2H���1[%�����}�KT+�\��b*��M	5�n��譔���f��Cy�{?v���Ԕ1ѐ�n��"ﶲ^�`@Զ_i�c��4l�67o���e��I�X��Xg�7�u��m�\���	�����J*�^a�=�X�$b7S�B�)+�Q}�)6���n�d6���e_78�	;��C�m��Y9H{��Zw����̲�T��cK�C
��;��R�x#1�`��X���o<��A��������,e|�{<�>?��+̍x�>������z�"��F� e�/qN*Jy����k�4�c���g�B!��>ۖ��VQ��*�'i����[9���{��h��d��6F�5(�IN�X�*�o���.�f{��Y�e�Q��m�����u��p��N�m����WO���U�4��K�
��gt��J��:Vե�����=)L���>+4(ZT�GOV{ W]�2�4m�dN�!�4�����?M���t���ɒ��AŞ���=���sIZ��ܧ����qd�r�Ӹ �)�"��8��n�=nV�2 �� 
�zچ9"��@�� h$�\񳄊��9&�)�РL9ߟ� ��}v��D���z�ؽ[<�zk�.7[����%�b��
��㇊=u�ٹ���M�wG������WM���5��f`E�� ��$�MO��=�0�-�2��_z�Y�("�29��U����~c�Zu�J�����DQ�n�5{G�I���1 �X�2�1~K�î��14���>�E:�v�IO�1c�c���RϽ����!-`mu�۸>��$�MZb���}��<�Z��e��\��v]nԗ���3��q�;�FI����^GG�||��P�:�WI-�H��nظ:�PVf\s_|���_(K�Hc�����Б�A�-({�uGb�Df\���H`���T=����3�� R��剩b��T���K?�D���G�O�j�o�8��R�����T�а��s�(}�Y���[�㖤��)Ĥ��"r5Y[.@��M�ɸ��r�5a8�)�֧Y\�=J�G@L:���m��(}w[������E��Ĭ����]��b�%����bug��ܯ(����M�8^G�D��0��r �"�r�76I���W�0�����;�C����G�N��
{�l��B�����a	�}b� �V��4�G�<��h���䨀���p���%�����
	�HAz�ˇ�q��b���c��FJ7|�+��ӱ�"�\o�Yx(c,���Lu�Ѕ&�f���p�V�!s��E����o,����SJ�5��)J���3J���/�$v�Q�z�0XT�e!���>�72�8�4��V�d�-7��p�6�%���:�ؼ��o�y2�HpQ����P9��h�'�ֺԏs�궞>i�k��妬�]��Z�$�^�4a�};y[��ydkq� ����n�~�\�"d�3�_F�B4C��87�,��E�����á-k�{�ſ�}:/��t�j�/����*5)����ۀ"�~uMN-��������
���9���+�����g��q�P'5�~��;��EB|>W�c��������6���p�}������t)`���VC_��=�GAkSl͒�3O�5�44����!H����z`P���Z9�-_�[�u��R�+�d��9ޢ��f��*Q�dC�ၻK~� %�i��	y�~��W�V��d8s�ϟ�� ,!��|�$R'h����ܖ�҂E?�%m*Mr�I��pl1�]�jTq���ɯ�#Q�������H�#��[W�jh�X���������[@�
���m��ɩX;٫�<s����*�\�r>)J�
���&)/O�F�A�6x���Y'oAj�1�OJ���ـ�����l��N6�Z�1���(P�����^��=��ti�g�T�N�B(�6��l�����_$��
�,��4�qjl$�ƙ��v{$�ak`��"A�	q��/��-N�l�+���i�A@np�	o�^��`wsq�l#έj>�� F�<������������3����fd�BNjZ�fgY������|F�Mh�R�j�Փq�����|���_;�c7�'&N^�p������QayF��KM2�*N|,⍸ϋ���IX;�6��|^.�C:�[ڻ�����2�����g�^��w�w������qk���pC�ƃ��N�S(趏�ӑ�48�N�~��ǣ--mtuu�t�	d�GL��#1r�-�b�}c@t��$�5kO��u��:�%˺&���sL�YnZ�RG�3뵻ۼ�����8�x��[�ws���G���;*n0����+��A�ͪ���B^������,��]fY�|�<yl���*��&6�F/ �d�	��Ҋ(��RL;n�CB. �֛�ŷGF�E���M�fC�*��f�X��RX;ωhx��������8���S^ih����>_�N�{r�����dIK������HQz
���W9����bz64�ɔ�IT��ԑ�_���U���%s��T��$0s1���s�9��.n ������ԃ�Bݕ��h�����:x4ý�A-����ct��$sMG��G��$r2�X�����grB孚��j*l !!�O�s�"��b޽���ń&А���z��XK1�Ԍ����Z`Y�e�C|�wr�fͳq�������h�>'�YRA-�pKq^M]G�.�O*��ʾ�U�al���i(GeVP�~�n�~O-�YZ(?g��Y���-A��~O�n�U����f�2�p0~Y��ш���(X�v�F�E;���P91D��Xb�y��um��G_���㹤ƺ���j$�&>6��0���2�D�.j��4R�8�\w�q��Fݓ�ѾKz�d,�,�S�����t/c� �v�����o��<(f�}�����U�JIk��M����&�2����j��o)�y���g�#o���19?;�������Xܒ�5��T4+��S��+�,C��˩������;7??3�[����y���3�G&s��9g<��KP��lWe/$C�L���j�T��L2��K`҆���Z�7���F��w������py��92�">��«:Ԍs���%\��������a���FEw29aj�ԹL�7;�fǷ����?�9��3ӗBČL@�~yD�0KJ��)<�;Q�=���z���@�P���������l$C� �{�6����lzF�A)�O6������C4����ʸOBA����b1��`��Q�.徼
p}~��@�@4l���[������&#��`�#aW�U�#��������D��b���&�hj_�d4�z�7�� g��{���0�e�O6��#���cP��$̫���I�\���7��[�K�19�32�ن�boQ������}�[ZT�G/�ԇu�=�NV��Z����-�Қ�$��j��?���I�n��j|�m����`A)<���aJ�a3�q�
�S�X���W<��ϗ|��F �%j����Z)��
�w�W"�/u��뇮����k�L��'�S�u�(�?�K*r�*��3�J�;`Fh&e��s,���f��sBt�A�b�W0<yS�'�^�������(r��}�}"	(bb�9�G�p���Ux3��~28-D�@��`b:�S�I��V��͜q@.�<�z�Bɾj)�儗��Y�^8�~���S+[^���o'����k�	�@
 ���X[ o��c��=�YW㗟��<o樂����r���Ug������,kh�w���w������!S\�)��(�v�&h�hں�8ggb,�%��-���J����<�Bbj��ޭ���?��K����\�C����f
[�I���!C��~hV�V��}��|ڊ�:�o��oz��-Ջ(���Ԙ�лC���>ژK{����0k╫��\��k�"5-�~Q��+��]��[f ��_=���x&g�d*6�^�9B��i�'o�P��K��Sܟ�>8���t��a�VZ.uQ�i�����w$�e�Ǚ/����:�x��y��($�Ws7Q���`j$D8��H�?�ɮ5-��ƾ|F��L��djD9��V�\%1P؅8���B"�I��ɹ�����[�G?L����=���I�4�80׺o�� 򖒫�h���+��b-5c5F�(�_�E���A�.C:��煹u���AɤA��k'��&sH<N�Z����J���,��C�NJ�"t�;Ԙ�|�/	γWpB:�v!�?��hk<y��7ΐ_��Uӓ��sqh�ѱ�ɩ�C��}�m����i�u�@�w6�(�w�'�k�$̸o��rKp)⿢&�}I�����H�x3 ��&��(��,�>S�:��t�e̅��'����''��r�Sq�-̫�K��煆?����|9/^z�#ʿ��yb#[ b�ت�xN�d37-\Όk{��^���1gӹ,����8+�>�y<Ǿ	hp��%ZB6%�E��\� �����j���{Z �8&Z���d�$UeR��1�o.�.����M���6��NN�>��9���|�����Ԙ��� �Ff'K7����t�����'7�������{�k~Id�2� N�qR��/���g�bȜ���A��(W��Ҽq�WFד^��[��d_D��kx9f_M�����LH�c��M�j�v;�p��?����q���a>�����9��i�9��ߒ�P-2o�v�V�����V�X�](�o�w�����Dbڞ,n:vV�7���˫!�_��?�2hք?J{�	���%��fE)d8��-�������[�����+N ��La­���@x�8�e�.v����þ�:ԋ� �yRY%���d��H$;�ݜl�t��)󮆨�:��bi�{��Nc������;�'��Ѷ��o1i�""�$��[��_�:s-� h�NA���Q�Ի-�z8���,��ST
�D���(D�l�7���"��X� �<�¦�I�!��O�Ǥ����N��Q��pu4���6T(3����t�I ����(I7e>-���&؀���Yy����& ��I�2R�%�0�Q�q�7��s�ij&Ih����Ss| s���FU�F�@��qߵ�h�t����|l�ΫТ'�B܄����o���3J71ͷ���z�אg��W�c���^,p�Կc,I>�e!#e���ⴔD^D-S���w�4�)�q�������7��{��<���<b��ҍd�{B��_�\�FE�swv �^��U;.�X2�VZ��N�5ל�U�w'���b�p�e DK�v�/�@��{#�Z�l)be�1�!��0f�z�70�Y5�/rd�ɨn09�t��M��p�!Y�a�b�P�roK������B��1���Ƕ$
�m����L��%r�©s��G5����(7?p��eWT���W)�|���%���.ߚ�R����#]�Ad�Y������SQi�h�f.�(!�L諌��٫����|ݗ����t�C�;TZ�^ꖦ�'��*��0�y�%�d�86X��c]�g�G[�t����-s���=�qp�&o�0H�`����~��;�UM% D�Dݷv.͹Ωω��,R�	X}�M?�]�-���h@=��i�¬UQ��s:�U���"�?Q7��� 
+�� ��Uhm}��v�Ǡ����,:;�(��0�H��(��K8��aWK��<~^�}b�q��q�ޙt���X���2%/���潴�ơ���~�q�n�؍n�؆�F<t�/L�8:��iC���F
����GDri�R��D�G��kǽkG}[g`���a��8b,`�٧�������ϔ�����K�J}kvU��ed!K�q����_� �˾�F�v~3;�Ot�[�vK�`@��sw�U�렷��+�����'�#Nxj�AB�"�Ϙ�}&����|��5��ɽ����98#�`�������QQo��0H*
RR��tw�(Jw�t7� H# �tw7�%]C�0��3x������k�k�s�ٯ���]�,G���쭨��GS�T�;K�/KT/��b8Uj����[�/���Fu����)���3�^�{���� z�g�fgk<x��%f;{w
;-���\!=/4㙐���/D+� J�	������y�ܪ�b�`1M5�M��z��0��j���b�h�Z&��8�E͞o�R.��_�Q���<���,=_E[ʋFr��A��F������2f�zǗ�}Gn�ME������mN*g�y��4r}i`�a*P�������8�9fT���4����;)�O��gM6��{��ƠDΆ�B����-� �ޛ��A\x�5"� ��(7����<Wt�Q��z�J�g�/0Ihpz:��ΛX�k�<��8�-�MRV����0����}��
�֒R�>�v|�>�o�'ʯ��E��&x�h��*\�n^����?��>*Fm��q���}e��&]�U�h���h�֨_���+f���ɬ���ᐘ-�� ��>�����<�6�c�$Q�7s�ʁ)>&;��XP]��
S��A���Y� Kl�2���D�-_���^���u2�E��Q����;���L��B�kv��ң��-��n{��o,����� ���cR��O-g[��b$�UpШ\���RE%97Y��n�A�$^�����v�y���PU�W��^��<ݢ�Se�]�!��ϯ�R}��$=$@���y���V�0iv�����Bv��O�@3�ϧx��2v�ï3�<�Q����)�/�e_��vĿ�C5ek\;~1�=�Ի3?!L���>�z�c�ƭ�N���C�|�!^�Ȏe��������L���<)�?��AX՜���`����.����~ZrrV'F��s��}8SQ
h<�gX�1H6��d!O(1���_93����֒�������\-6�̛����`�,�L[?��G�b�X86n����p��CɆO����o�Ǯ����m��+Q�왹�C���b�U<���8��QI������:o+ݾk@Ktk��7�GƘ���nX���H�����nl!{����_sFN�?9���<&Z)��枅Bణ|�T\5xk&�f�h5{8q�I���Q��y�[f�w6�E즊�[���h���:�X�)�x璏/�@��A8�>'?��=��baDC�@����]j�i��
�(fz��x#�D�/췾�{�߸5�N|{ �5��Δt���n�C�a�/��15�R�7Z�A:�E� {�ف�������_���O�reK���6�a)�V΀'[��[
����P�cF�fi����2��3��.�V�mX�P��vڌ���Ǖ�u����sv�E˕~��	Q?.�ÑYc��3(3d����#3���t=>����pw{� e��<;�a� ��G׉mu�{��R���T�b-qjʃ�"KO�����荖ġ'��e)�v�!z�W�(�K$���yf�������i���f!��h|AQ���%�Q=]�;��
�����6���G%���ڡ�ȵ�T�T��;:��|J�},���yi�C4��H��g�r�����I��f��N�w?ʕ���E�� 1Ǳʦl,������S�%�gul#�[��ߝ����(�&�ïn��Ǡ)ʦM�n���8�O����oN��=��ohy{�"Y��Q+��C%���**5665���i�T(/��k
���qx�ִ�������I�r(��"$X�p�#ZZ��'osY�z<!��>Y>��O���~n�Bt�F\�२��m���Ub��� G��B�5�}����{�>ewX��?�n9O��LI�)��abJx��l_\��qSūȖW���H߼x�����u��e��G���Ⱦʜ�Rٶ!�X���V�6<�`��za�;�p�6�e�;�ͮ�~�Θ�m�na!RE��~:���~& <Q�'%Zsp�����EN)X�~8����"�+���SB�bl�)(�aW����R[�<#e���,-d�|��$X��=����� ���u���ۨ�,��$$�A���ɶ��s����2��d�tcr$������b����[�I�xʜB��KQ�z}7g���{ro�r��sx��rML�n�2��r$;���_�Ơ���V�iz�2Z�B�����r6O�]���A���k��M���m���}�_^-���5�x>	B[K����7� g*�v����:�ݚ�@�T��!�q��i�<;�^{�8y�I�4>2�������cy��mp�[PȺq&����6�֧I���|�Q�����k_/���#d6ex<�}n�~���=�C~|�����oj���=�.>�,A[���J�mA ��FA὆���!���3�����P�w��Ǜ��uL,�u���FM�g��R�@O2��f 6!>�\��������} ��Ge�c�b�c��^�8����뫇��������V��h�w�=a���*���$B��Щ���!����
"�$��]Ku��9�=�uY��1

ҟHc���+^��b)\b9�0|��h2[��+�<��c�uy�kBrOܽ��ѹ暰�}�8���������gm֨#��B�@�ڄl��NF3�E�D�<WY񽆃�M�á{fV�	�Mq˔X֢=��s9��gκY
_��"�^�k.�� hjڿ �N�L�/�3��Eߏ.t�{OL~�hYiٴ�Bg���NN�*�S�U�I��s������\�c�Ko_��A�^�})bD�������!�%��|�ۦr���H�D�tdB�����f^��!"[@Ck
�)i�rx��
�������A+E��/�k��u��Л���>����T�|��/,x��Ί*����>�%��/;΄Ҟ�����9&��:>�W!f9�_)U���2^v�$_���7�T�r%������\�n����l
�#\N�݄�A݋p���R�>ȹ�O2c�etͭ���I�(죥�iAg���T3�~�5y�^�gj��
RB~xʥ��nN;�t�s��c�|��u\"��;j=�{M}!�=Fpw6
��R ���ԉ�T4�}5?D��I1�|$�aV���˯ۅX����6b�D�T���%����<���֤k�*��һ��6:��*�ߕw�|�06᝕c�)��I;k���GG����fm������+�S�/p��x�=���*��������s��2���y��w�:t� 8�4u���-6y��8������`&�b΢Id0��W�v���&���9e�!N� ��r8Bjq���
�|�
n>bn߆l�;��|ҜG��1}#չ��"�R�N�����X��iTI�5��Ю#=��zY�P��hd���E���qrA�R�Ş{Z�,��B5�b�����6TެTN����U��A�9���4�t��~��)y� ��pX�h�}+C�_pJiT�W��)�����(�>��r���<��0?M���oR��S�v#��%m���1_쯦m�4���{��t?�i��>��}Ʋ8�C��g�V��J3�r5���[�g�:P@��҂�#L�{�ߖ���Q���jQC>���|;�>�a *��Aϋ�k�ю3҉��B�^қ�Q�[�I^��c�7���;����88^%U�2o� 
�8>L��R��S4����:�O�^%]��@g3x����I�����K-{�2�}�޵ČyW�_�����Ϧ���!��.���2�(�=(\i�.댡����t9��M񜐋�s��h�O���=�s*�: }r����}��r\�IJ*S�=��)�O�/'��նN�$?�6$��Ъ�ka=�j�Z���Yٳ�PKdb�5g�Ma�f�?�KɝY�+�7��'�R� ǰ{~=��|A�{�����m1ɃC����8-�������..�ǡw�/f̻�i����z��!������R����J/]
��9W<�BX�� )�����ϴ/ �{�1%�.��9���RPg�K=��o�Y�%����éu�bj��{m3�p���D�r�7�!�٫ �㶴~�sþ4/u�4�ȯ����7p�]Bͦ��~�����-3vcش�b��~����␿w��!&z ���I�C|j�ϭ~�"�2V��%����|�C8|�ߪ�%�V+�{̇����.�⛝.Y��L���r�%7�:��L_
��ܛ-X����!A3��/�q3Z8s�����lS���k�N(1� �?O��G��**�-��k�����ԍȧO����َ&�mzcd�A��Uy7��i���Ϧ��%.��� sÈ̔�GVe��Qc�lFcp�ZޅC8��=�^\�y�)R�q��}W����l����`�x{�O��A���Ū���C�'~�eA�Q3������3E�ܞY^�`6��9�8:r��C�ʗu�|-x�����,JV_�c���?�E�I�>4�P�2d�����1t��i�4��t*�����3�ir����R��ߤŔU^�m��b��x�az��~��|)=��iua�h���������GQ���=���ݺ�ӗ�G�ĺY��t���W<ٙ�46@<�v=�M���i��&��C��jE��+��a׶���L�=n�G:�K����`���D�%i�i � �ݎ�����]�m��Z%�&��?�P ݨ�<V�.3𻪍T��
�UGDO�I�3�w�8ke鿈�&��0�'��B�n>J�U��0�� \b�R���ޜXXp�����ˌ�Y�:7��__P�{'��&�^e��?%-�'
=��-s\�#�t�����T��0����M�(2s^�E���#{:p���(�.�fx���_dW	~��.=��t�xb26�� i�C)�F��Ʊ���W��L��D�n@/X]E4��M��]��]�r�="��>x�;J�xgWv��~Y��Nfs��qé���J���f��1]�����q�]���x����c���TD�F��$!J0�Oth_�U|~v����7h;l�-3��������?s����ꉤN���="%u�h�sڜ2!#J.�C����v���E���������?^.�Ru�������w�ޣ����8^iAgy=�4u���:��)�^E�����F���7��UɃ��>Ծ.#a�x��+�͖d���Z���A|<q�ا�}��4J�����ƳO�O�+2��'�*ȟ�@�S=WBټ����d5�Q�����]7V0z-�d^�-To�u1�s��)��j��Q[U����J���K?�L�&mX7����U3ݗ����^�Q{�0��>Ԛi��
<[k c�n�3 �?��Z�~U����,b���`�  �5�����i��c>���H�:�I������ �zA������-�9���8�ܤ\u3/ȃQQ(ް=f�k�g�Ph����wL���-�O���x��V��=�s�?�&A�E�D�c4����m~�.D�@-�+&v�C����@���f��BL��~�gQ��A�FW�O�%km�쟴�~1I�BHE��#kD75�k��+/�L���P�վ|넀Y��=F���<+�p���>�c�K�-�	wz��[���e��$TM��	�<!
���~����ð�J���4�4�E7Vb�}�y%��T�M.S":�A�= bߢ~�q�X�H�K�_-�@�Ь���r�!���ׇ^����E�/���D����<#��-�&�Ov�P��^Lf���-ˣ���>�A��&�sg���v���íL/v_��~��zi�gH���Stk�B�����d��Q4��ۗ���iQ3���D0��I��a�M�9Զ7FC�j�5�!c-�J�l��=s1MoT��.{��5;C�L�y==�*�c���qk���"g�zme�㢨�ǚ�=8��!�bw:n�;P����ʥD�@�}�w��ᑋ�m&�	:33.j����V:�q���&�^K�|E���S>��3�+`��szc��B]�Z��q֜�d���eMH�{�����)�a���Q~����yғ�����r��Eɹ�'7�ͮ�,c�	p�$���A��"�b���>��2�}�n����?6Q��%V���-��ȥ��7\à�?��ar����	?j�p��*�FO�ku������Eo����)x���Ý�h΍��7o��I_��Z��Q�E�t�RLzTpN����qfv渰z8I������dZ;qֹ�.y7��"�	�'Щ�,[���J-^�`2�_�G�իX�����Gq���VG��j����
��[�A����7�6����䂉=j�4��Fj�����5q�Z�	�|�����+�|�g�b��7���j��Z�?:6>��� 7����\';.��T��$�v�.���;�Kb�G?}<��$���AaD����=��gp9�� �����p�N=��gZ�����ɭ%���'.��P�qdF���7���go;��0f�3��_��hs����m33,rfWE�}I��C&ʴ�S�
 ��<��_���H���u��{���:��L�'�MtZ�����}�^{y��R�����>6�8ڐY��j��P��*.�&	1��L/�$&vGW9|C �mec4�ె���,��u�Ǝ5<h�3�c�}�| �g'��\#�}*�#s�?�bbKK>A�]�2z*�r��쿻��G��Z؉�m����j�|��D��"�?�������keƧ+f� #��\���A˧�R�]b�zh�uu���}��g�ߥto�Q��~=�lx�q]v�?��1o#w����f�R�N������[�>������5w��ιQ5��*I��0>0i�C��Q�~�n:����BA�t�NSH�����>!Y�G���e�[�O��J*+Y>����4��OE����>�9W��f0����؛*X�����	]/��U���ЩR�*�Y�1 ��c5Wze�±����u��-��ז[|�G��n�^�;Az}�D�)oR;S3z8�lAJ?.E��Η ~�ߋZ������?�r&�dO���M�d�2t���uń��svqA�#T|�u�}��p8u�π"��-a���J��WM��+�`��sX�g�X�]��bs��� %��^�lZJ��!��m�|��}�ި?�j������.�B�As7PTз�<�oZp������i����@�.�,��-�����ar*Q\����;_v%���hFBRbS�u��u:��,r����,dF�֙��\i����M�fK�xp#L=?6���n[q[A"�?io�F_CV�W��@������h	�)	,��\���n��4]��#�^��b��ܘ�~Al�B ]`o��/?��\>�e?���Ln����|WQ�ψ���_� ��.W�k��3�?�*��q���\-KH��?�R�f�Z�2���9\Zy�ji��c�RcI��D���J'n�y-v�Z^�[L�����2�qӅ>='��(���bQ��̄�����g�T�{���d�"�ϡ�tK��)���T�f؁��'�9rT�QL�M������7�j�%/�Ÿ0"���v�Q����ϸ���i)��I6吉����y��+/���=�f7��G�ms�+��~�I�
��t��(C���3g��w�i��j*�hӻ?M�����^o��K-8���{��?�lG<ɿ���x8t�S����ɻ��P{M�"vo0r5n���[���$������]�P]ئZg9�o��޾��o��w���w��wl���C®菨���dE�C����M)���0�����M*�-���f��4;��C�[�S�2U��I��q��ɚq�����9V�;Nq��Dn�:��XG7�Q��ώ�Y�q%���߿Z����Y��0`�W���b5�h�K?�� �^hDts�V��č�-H��(��pZ����f�E�<cU����t�=��j�Xk+��ۙ��Mv��<�V]�	��A�9s���iG'�3c��u��o^�{�>�ԱE��1�K�t[�{�N�C�MTi_m����%e�RK-�ۀ��gm�QpJv�ģ�?:�:����3�VZhQ|���|;#���E+�c�.UZ��ڗkX���ل'��9���=Ѣ���j��~���r�M}�ᯔ�ԫ�NX��XYֽkiD3�����}�⠧4��~�H�q���d��=1����cxsP�Q��O��f�9J���l�U"�!)b�/�y�@��T�'Xz�^2��¸�������e}��R"sOP�� p���0�1�|���n�~|��uVR��
�����7V�̂F܍� q$.�Bqۨm}2���\��������'��v�����Zm�☒sμf'}J�FOkhH�l�V�RA�.�A[W�赒'_��}}����K�&%��l�غb7��Q7Au��L����obR"$���G�޼����3�j��c��?H�}:3u�����= |����I�[Q�L����b+[0F��fA���.v��r𔁁��%����,�y��?�h7K�T�s�7���k
�V���.s�1y��X��6�$����4w���q�}��jpP�G���g���o��ju��',h69��BڀzuǜԄ@I~8��6��k?L�Gu;������~Tm�z����� (�u��³��u"_�E�toX��V��qօ��	�p���J{na�e����:��y�n&&~��΍(���y�E2G����L�O6Վ�j�U<�%�Z�y�ǜ��=h��ocdo�%o�*��dR����ZI�c�q]o>m%�"�(n��r+��'����G��_la��#Y^��9�Y���b�<*]l���`�I-�y��*�� Q�����Y�`�y�5��/m�>�3p$Z�s8$��6�^�'BϚhQ�z��c��k��'L�E�8~�Y Le���vUe��q�J�4s��i ʔ��d/(�;�a�ըRm���-��X�x�a��!���i<:[��S���L��VN��3]:>��?�o�����e3s��Q�غ6�4�RVݤEjG��tV�@~� xr�޵j2��h~_[W�c��8er&!.���2��U��V���[� �J]x$���/[�~w�.}�|*<���Z�n��t�B;�jK<��~����pU3�Ԁ�h��,�`��@捞��U>b�[��𷢕��D�%�ͨ���V�Y�7]�1O9��ku����Y�I�U�������[,)/�ٽ�����S��1�\�ۭ�B۶�g�\&��MCS�i��P���/��J�l?��uB�ś�ɠ�q������R5*N����ن�
9���⁑�}Q��k����k����a��CNĊU~1|K�]�Y|o���v�t��#;��9��RGu�Im&N�f��f�b����Ë������j�|;o_V�T�����S��w˯&2dOoN/�e8�ڻz;V��K��,��x��S	�w�G����6}��&ː�j�V�>@���	�����f���3��Dn�>��q`�Q��o��M�{��xn�mx�I�zA�/�4�+�=��J�)����q��P���,�/2~��e���w�P`ՙ5q��iz���+σFɜQ�'g�����PmX���,�213G�J�V�Pӡ��uP�*9i��ۯ���nW��+��珧�Uj1P�C-��t���y)h��J�&���J���E���
4���oy���	vU[��'�|����16�w���K�ꐨ�_O�����/�9��7�f_��T��-�=ۡ�-��g�h[*�kG5�g���Ἑ�)��81��c(K� ������|q��7�W�  �N��u����$�;��v�kߜXX(�F�j�۝R��>������́7Y'{�`[��烝�S�w��$ܟ�D�h
��m٢���/��T�V���`�(fY�z�:پ|��<]}|`*��q��.ߗ�e�41�cj�:�����6]��]dF�}:��J/:#Ir�n�~�joSP�}�e��nrͽ�����a䞁0�����<P�s�(�ЁcDI�vMѨ�gg�Ǉs��K�HrO��Z�ϗ����)���i�C'�AY�d���w����b�����x`P�PQx�9C�S,E�!�%���k���7O��ށup��q�A��̼��[C<u���t.#��<i���]!��;Ī�<W�<*Z�WM�������(��k=�C<���؜����q�;��g���䖉��a8��0��5!��U ����Q$^_��#���θ�ضk�hWK}h�@F8-���n�[�:U��u�:�'�!�(��=�/�GEpӅ��[W��k�oH2>R��NH�K�f��^�Q��+]�����4��Ex�Ŝ�FU�"�!S9� OǾݼ��˒�X'PL��h�ә=��}�I���J��}IV���E�+1�K����e�������W��:k��m��}�C�A�ڃ�h�ͼDD�����\�BXB��W_:�=3�;r��pV�4I���,��N�!^�f��L	_V�o���T�<��2�w$���D�zhZ�j7۪�ZɎ����/5���#�.�<{?hG���5U#FĹm}�A��8���1:���%��F����\��������Df�+0��	ۯ��
(*k��Az��+��ɾO�{��A�J������rm�����=��l���@qFy5^@�����2���Q4�G����OBV�6��1����.���f�ޏ�p����P<.py�'�!XT;]2g�ydܾfbR;w����ی�1��a����2�&��<��<)^]�x��#�A�%���e�{��Z�.��*{��(Ĭ1�ݩ� ��	x'�9�HS�i��.Ȩ�m��t<����5������5�,�����������U�G��Y�ߢEYW�k���o1�Q���c#ѺO�4"3D�CA�C��{Ϋ���cs��8�,��+�^~q>3_�lu��>�ti2ZbKF��Ny��T˗*������: �W4S��|��τ9���4��l%�u��/�k>	�ޅ9��*((TQ7�pq�)���]n<�P�PM��&I|���C�d#G7���DN���BIPЀ��V��N?ٚ-�w��l���!T�	�{',�{3����2��
]��V[�/N�އty�-�A�bѸ6u!tJz��GM.�PLibx�z(�����yL v������|@f���m��&���7{@xw}�aYȈ"ȉ�i!��"�R��F�k6�4l
�%W�d[�
����cP6	����v:�MW�.3e�P��)xq�q�cRrt�{�-�tm-j��Ւ:C���V_��σ/�G�%��D 3���vt�
�n΁��/:?����Hy����:Z�ǹ�E
���Pm��l�-�Ow+�ATRK�D�MB�r�>Z\+�϶��`�)zsC> h��nıyH��ep�ݾ7��go#���������L�ؑc��ҧ�l�@
��ړxX?�vֶ�H��~�0�%9o���.ik���a�Tӭ�GW��1 M�}�%�QJ»^~�ϭ,�*�ww�Vc^����̸>�ό�X�d�t�M��h�wP�CY0�Xj�9kC޲��	�(�PG{& $!͆�t(�ᗚ�]��bF��ug2s�!��A|OM�$�<�K_v���=�x�]]�@e���'E��#tj�dÄ�(��."����`����Q��)������h�J��ͳW��w� �+!���ڌF|�$���K,PZ�l�y���`��d�zۆ�u��5~��|�M�������L�Ł��b�Y�r9�t���,c�Q���y����������hM��[�r)Ϙ/�	�|�-�e  t�a �Ybx:]IQ�`��GL�VWUwαS��s�ï�^bO9J?��2��m�-a�=��t��:Z�[a���wF$�[�K�y)/�:Bg�6n+���V�ޛݔ��;�1��d��(f��"����uk��n8�;y���@>�]�w�����8���}@�kH��68W�ڟ4����ͫ�q�w��#{��(��}�������M~Pߵ-�i)��}��x��������0�X�n���1&�\��m��*m(9��B�3��S2��(B��>L+��p�)�B��O�Y��m/���Aw=�	.��j�B�?f?�n��EV�{�k���N�^lx�Iq%vF��G0��J�ĺl%@P0�1�cԏ�d~�S��F$a�ij
T�5�cj��z-\=�� q�y�8-�+m�cLk�]�}�j��sf��D9��+�#������4����yX���㳧u@7v#�b;:@�>�����[�!7+s�X�+z<�jX=Ȍ�H������0�C_�:�M&�?����1�-'#��ǲS���N/I����F#ZJ�U�8�:?��&��y�R�����S�e-�������j�$��]��UW��ҡ�O��bZd2c&^�J�0B5�o�| ��b�S��f{g���h�3��	`汍��2�}捚�Yq�����3q7�R��u�ڍ7�` �������.'M���.��C��k��Q#e�},��a|�XX�S9H��:E�r��0碉�ĵ�_�㰣��%�������|�7ʯFs݊�0�Qz�6�nk$3�ü��w-�>bT<�>��4C����]zZ�ۧ�dT�$h�����ȗj�\�TD�0��w��>4�\�d��<�2�L��k]@���I�ŀ9k55�h�X��2��{�z�)��ԃ-������b�2'e�`*X���56�:,f�+�Nn���'���6F�M�9���^X�~�㛤MuS�P�ml���c�LM>�k�5 ��G�w�Ʌ�#H�C"��[y��S�7�G�5R=�J��d�::1���MtТ����RT�g��`�y+~���A��탣��J7��a߆5���}\{��&��"W��c�v��άO�=�>�����^y�0�.Sf@)U;�C�W�ۼ��U�ˮ�Ȗ�8��D�/ze�S��
��[�����.79�5��dJ�>���$>g[�
۸�"�i�^﯇=/�'��ù�/ݼ��%.�9��ʭ "�0��B���;�U��Ŵ��~�� ���mM���4gJ��s٩[iIK���Va���+u%"��/����X[,l`�2û�'N��X�W�l�f|QU�x����]���U��_ox+l�Bk�o�|��ؘ���X�� ����DMzvi:Qy��Cl�#Ӌ��:��݇��e"L�W޺�c�tP��mW<�	2�Piɤ�5���
%�p��޸l?ýC�8�T�9jbQ$�-���L��)Ж�����i�j�M�0��KĤ��<?�z��C)iYY�x�w�ثȶ:�̱���j$�jn@D��Q�% ��G�!�tu2�����qa��/�t�چ��+��-^Ξ�~�y�������"��!\<�!N
�R7��*�f�����(XN[���?��6���9�
Pt�'r��+
�0&�*������fc�DV.KU1����p��(rb�H��g4��~�՚�1qr+�UDk~I��W<6q�==�Ƙ'�w��N���HE��S�+�G���F<_P���.� �}�~e�׉Q-6i_�K�h����?�BZ=bب�D�%������H
HϔIx3|/*�������禆�_��n߇��jX������,gŨtQy���!������3��"n|� ��5W�,�[�X�B�ua�ɞ�+����4�� �t��B��h?!�n��J�Fş����4���ѹ�XA�v�C��5#F�Y���U"��n��~�\��l�L/UB�%U1�-�|X�L�\��}��WQzTI������,+�/[]V������*��L�'A��_v᤹\D��yE?�7�6ͱ}v�5��eN�M3P�-y�*���/��x��d,x�<�2���y�c���^Fd\l�I�~Q���5�D(�C�[j��n�J^a���������#�/r� �������=��E��9^��(�If�ӕf���Ȭ�Ui�Z&O��YS�y*3�tp�U�h��M>��u�kN�����3�Kg�3/�\>F�J�i{o������t�x:�I]���6Az���ht���mҏ����ќ��iV<缺��e���9J`]�٢b���|y-�$��zk(u`�cW-�̥w	�I�im���ʷ� �w��ٹ�Ɖ�׮���+W�j[( �=����Uk�T-�x.�[="���kD')���fX�Ie�2^pWU�$	�n��#�Z�3D�a���~�P�0_�$ �fml�|��躗��O}�f�T��A����>�B�*����5�S��E�a�6F$h�'-~?0����������op/��M�_�=���3#W��h�kiC����4^]���.��ީ�\:�Z���I�F��S:��`4�ii����t}ڦ���J�BXm���rW�&��\L�R�=޵�`�,.l]����rwO	|��[�N ���mm{���M.-g0wh��6�u�W��9���BĈט�>����'��©���u#�ENr��x��D_мk
��w�s����Eu�҆����j�O��u�w'���T�����#]���9�F��K�0�fW�J��,~z���U3]�X�h���R]w'9c�~=�PV��a�U4M�it��;A��D�����a�&��:9�MY1RK��72�����w`O�-��S���6�jW$��[)��k=b��նl�	�S^����K�p��������
h��5��>k�5y��J�������@�oPå,��^s�U"�-vS��[ȥ����tn����J�-S��͟|h���:Z�zI9�?FBGyӲo�� a�ԟ(4~�;�����������T���q�L|D����v�������Y"}���;�Y>�l�?;�+tH�i�'y�{3�����i;&��ǎ�4ƞ	)�
�75���0��٫�����Aץ�>���8~>"X0u�b���y�@�kEK��ț1�o���$���a�w��*�SmH�{�aR�}a�x����N���J�3�����x��c����#�`��L�mbvк^�{qʁ���0_Nm�����v�����qz��n���+��a�_{�Ոh�6�ș{׸��n�+�*�ɚ=���( H�?�ٽ��x֖D�& P鳝����@�8����h�R�eX��F^���!]�6�o^׏���QN�� d$z�������Fs#새�[��/P(��Ur۠�r��Լ�-n`;�nT����5�l:Z��-$�r9���!��qd���m�-	�ċ�~�ې�h^��n��,��V�.e��u~S����{�?y,s�ǘ^�ҏ�{/_V�W����;h�	"4�*Q׭3�o��r�iX��*G�,;$T�깥�Ǌԩ�V2���M�:`h��S�M>
M�>˷�;�(��t3H�z�A�/X"��m�E��!g����D�g�z����˚�#v��M�J�V%iڐ��vo��Y~�z,xS�9�nq����������\��{����������X_i�u��)�{�Ķ`A������~Ƌ�t�34q?Uru3��������އxc�������ll!���m-gJ�)x��k4O�7I�ޘ-�ښ��t"G-H>�s�[�֨��h��l�jM���ٵ t�����{�+��������I:U��((xT�-\(Ɏ1ł�b 6���Q��Qm���)1V������F�g%�w =��1_y5��"7�K#kgvR��<��]*v t/edP�$�w�f�o4u�|O6a�bg`�K��=o��Kr-�n	�o��'��£��ڞ��8a���^MY�����	@�v���ť򱓇��Ӑ�Gzd�̲��:o��m/�KP���ָ�l��ة˫Ku{ו"2�{�Y�v��L-��Ĺ85v]4�^[�xe=���S��HOm��%fP��5C�ʚ�m�����g���K�/N�
�C��a�t��o�i��E�K?�M�c�:c����k'������U�.����˂�Q.�؉Tۓ�kc��Cը�[�`�w���D�<�9
܀�Wq�u�81F�Vv��EGv���\��i��#������Fo�c���yĮ�^ �~�o�<͉]z�/��cE���t�(������o瓹�o�.S�'Ma>mML~������y�5v�.N�a����]�UM}_��đ|�_|i/��1��u	��-B;Aq�E��B-nA=l�{E~�~��|�#i.��<#�4�����U�C��`蚙@K7�ܪ���i��V-~�0מΨ�R��-QI��%���ΥPtf��{{oj���$��e��� a4����8MSM�|$�ɾ��~�Vw��8�����c����p��0�42�/1g����n���j�3MGD毺�+m��柭��xl\m��g�#���*s���n�zZ��e��̕��ޯep���GRڒ���5>L�˸�[��ߗ(��U����x�p4��[B�(L}@�}r�|C��[w ��]�˶[O�ƽS���:Q��m����/~�k2��sp�����x�{�7�;�es{M��j�:�sw�/��T�P+����1韜��O=E�c)��m£Y� Je1ZX��@�m6����Nk������^s��I)d?q����*�N���.��gҪ��O݃/���CBU_ yF�����{�?��e�.$h�YӰ�}����km�y�W�	��9��i�Y�S��<{�3B��^Ǝ�Ӳ�g_�����"|�_V���͵E��v*�^?�Oև�8D�Z�T��]!f�2�Ke���?3L�@F	��սr}����\ؤ �e1/ �[oW�u�!�4���Bp���A���,����K�{������������t�[���}���8˴F�E~/+k����J@�r�i�,H�Ϻj�i#��[�D`�װY��nCP�"X��z�?ލ�铖y;�������(Ƭ�;2�Q�8�+�I��;ln�M�����W]:�-&��M�� ��m�y�vT�Eϒ͠�|�<�:F1e�%��ѐw�~�:���^�^�[��;{�l>;���ԉ9�[�m��|��^տ�#����Y������0"S�R�C�����>R��-�&����mm��ޜj�{��Rl�vQ�h�j/=Qo����Q�$��숺�մ���b�,���"��O�Ά=nL�3���������x��g�7�$��O%Y!sqˎf�2�E�#9񜈚m�=R��_C3�a���H��*���v(ݫ��ݡ�
�q$}~Q���l��� ��
�&[�����ѻͯ�f|FYQ`.o"O���`}1m��#55���������'r,L�x�|^V2���N��$����xg��ʑoGv�[)�[?r1B7[��e�z՟�V<]1ؖ���	��c]Yi�"qt��I����l�B���i������:��T���ڸ�@��&�yt5R=+�;#D^N�v�f�׻L�L%n���l�ѯ�^����K�}S/_�[k�M�(8�GJ����)b9�3,�� ���͇Bx��[݅^�� z��ү	F���gđ��� �M˭�����&���"���a�pT�A��rå�zb��Y��^8�1�d��G�g�_�%e:���K�#�IYB@o�j�U��"{��%}�|�P!�7;uA7����~�7	3��=ڜ��&��G٪-"�����b��ί`�x	���:���q7���Fg��>`�h<W�&��� �r��J8�=$_������&���B��՜��:mt��!/?�(�ψ��?��J��n�w��"-�	rg�~IӥPg��j�(j����z�lQ 9�.���8%*k�i6�����ɯ���m@����b@��(_��$J�h�8'������.��ņ`��ˡ?h�[�b�u�?����K��TƵ�88���x-�}vJ0�(�9�D��]�_�<�1l�m��6@��k��*p���ld#c	�{�l�Sѐ�`Z������2�l���%н��;[�b\��r��+��Ml
U�C��n����i(Z=|3�YM(���-نE�CM�Ok����߅�z��G��m�C;,cE��&)q���i�"��*N���Z5m��@+6�єO�*�ޖH��L�v� @��W�l���</�֭��i�o�ϥb��iQ���%�gß!�N�#K�ݭhgS�)*� �?n^�8܊��y]���:��w���(��^H�(��	��Z/q�$!s�F�l��n���b�~����;����Sq�ʊ�p��'ea�+��D�)�]���������̴����(E�Blx�g�h�/>��AH��Z�����,��:�QP��Wi���^�����'�� ����O�k����R�v�������~F�'��=E�_�O�/F���k#Ͳj�]����Y�4�z؇��]��Ć� ���S���s�t�X����T�ߏ}=�蘙�;Bqn���o3�<䴕���T)�mۈu��mc�>riz5Cϗk�_��:c��AH��S��0�&/�p��o0V�;�y}}��q��1h��C����m�)����������T�W��l&�K�m�~��_ۥ��:6�_9����#2�bN	�U�j�B�vXOweݭ��.y�0�6�|KgeJwٍ=]�}	�������+�_Yb������C��m_aX�P79ܟ[�2d�3$k��>},gKм2�#g�=�j)g5[e��R_=�B��� ��}�%��z�`N�V�+�[r왃�ǷqW�%.F�w'?��I��U���?Xp�<�,�J{���PZQV_�=>��O�;o��qy8�����Po�P��cW;ԙ<���J�V>3^9��AZ�(����P��f�+�*S��%�.]"�6���WT9�ᑀ+b�k'O�k9Prj�G&L�4|@�D�D=�X������4���A �.�!<�O���Z��$�l3��A��(� ��Jr|�s�3�D�Ĳ&��[��t�wg��W!F�Fp@bj��������~�<�%�'��O���� xN��b�,���s	hd��yo��e�mCD�'�h8���rE$�/�RУL������2�]���2^�ڿM�� �����v�?�o �q��w��(X�EG+]�ב�
����"�g�}!F=�xd�<����]�!�JqM�����ۗ�]LČ��/	�q�5��R[Nf�:bd�e�J�k_
e�ɞ=�~����ڦ*ߺ��VF��:��}��/���+r�F�.Q &�����9�K�=H�}��rF�\W$����Z��F��
tV�^�;���o���'xK�."l�]_ ����
(Iߞ�\�4�����j�Ez�;;=�;K�����S�0V��]��Ik+J� G&Uk�ߋ{{c�}m��;+�gc^�q#�%��0����=����織,���]�t�i���m���BN-�����Wdg�"��g�?��	��\�B<R$�jKgdPMf	�8Z��2���2���xG�w;>�<�-騷�i1z��ໂ�0��;�N
��̲T�l:t�Uz���@�U����Hn������$xl�Zz&�L|ן���걛�K��H�[����|���o���u���|{fY�wv��ت��p��{O���N�J�b	��M,X_������y���_��<���ŀ�)N����f���_3�;�����$��>�u�8xxʭm^D�g��5������x�T
�~��\���'�^��x��������#B����jqD�c�٤kՐ���������,���_4���y��QVlA�y�gD]R>�,ȿ}��w��Qi��� ����� V<����}�K؜Ax����6|�=��Y���߃ES�S����35��i��}:��Ӏ�Ā辟bI��[5,�6���l~�tM4�r�U��� A@����CL����b�wA{z��i�k]��u#e�OL�sWg�\�h0�>�xn���!8���&:
�x����ϔ�7�m�r�7����=m큂�|r��cΕ���������x��U���rR�x>t��v�<��L�y�����r��(����(ܒ���XB�J�jq�z]��,R�|J�T�6iAC�������=l���6�V��=!�:�>5���v��P�r�+yb����^���n���F��V�A���n�5.G�����p���������x��	����
��|��qL�_���Mi�8g�f%�&^t��{q��GBN���q��9#�8��z�K&f+��?��cQ�֫�<q��_�ϿK���u�9���.,�w�m̗��T�P�Utӆ�܆�����60@�x@e�����X�_�������A��'v��|�d�k�ܼ?�=d�p��x��ʮ�nL/�9���"�֎��P ��ٺ�l`��Y�����~�p^�F��n�����l�5����;�>c�K99��d����AС�ī2�eC��}L-��	��8�}��*pg1f����#��·g/ߟ�^��[�r��<�^M�?��a��F�e�?*m�Z|�j3Oq�l�b� �W�2���^vH�_��b#��MxZ�Ѻ؊5$��;�r�,�T�w�50m/��[�i
�>\� G�\�
�o�K	�H�Z�֒|�
����-��,:P��U\xo�uk#��C	�oAe��a�(�a"Wa⣅�g&�l�g���܋������n��S�N��~�=�J^���$�^�mK�⡙<	�Qs�j}�\�J�@U��x+�� �E$ANE��Lx��=N����Q��x�f}q㠹����#���gf����z`�9���{��{�0�?��w*�~9[4�~[dt�����B��7�EaĬ��@b����:� �5���N� C�%���/}��V�M2���el�H�!n{�n�8��Y�$�H�~��7N��g�ح]��.��� �{`�d60<1۠?d���xv�}��HE�=k���o�� �cX���m�n���).������Q���t\�>��K�����g�|�{s��B���0���s�v�]wrO._o��.G~���&ƺtV�F��N`���d	��o�{*�e�[V��#7��a�q�~��j� �"����}��A�{����ˈ��+n≅��R� �N�]����A������u�͋TF`W6ؼ��4�����)�ʌ�y�N�CR���,�q��P�^����i��g�J�E�[�65M�,X�vfs%��� '�S��� ~�%�X����q��L+�߮��ǿi���T�䅑h�P ݃o}�ؾ?t���������^������tz=��TP����T������%ר��i���a�/���nbF���������9�0� �LQ_���o��"���"��WE秲�۞����yjl.������I�_s]q ���hQt�D*�AQ�f�PJ�D�b���g0X���͈��|�^ʻ�u��{�v�7�ѻ�ޓ���E~��j���/6Dro�tٸ4]��9����a�z�G��Ita�g:2j��?|m�Ƴ�-(�G�k��c��йrg��3��Kȓ�AZ���]�c}}��O�\��E�]��>�T�'FJ�Ai�A������GH�&s���+�j.G g.��a�����1���o߄h����j,��;
"����.rJLЀ0Ż��jיjl�=2oߙ��JCX�xM�`3��e����p�r�մ��i����'���&�]8�jV:��6ծ|�[��܊Hc��,7z@'��m;O{YE�"R�[� ��+��]�Tit�BM@O�!6ߺ![����kA7;%;���GMRA��Ko�d�f=�N$s�W��ǭ����+WA#	��`�fCk����ㇳ�`z�8܎��\���ux�1zĴM�D!�ߡ��c��?Y"�,�d�W��%w�ugu�*sd>����F��4���
N���B8�"G���e�#�f(�U�*�&����F�������-]�d��M�x��2�Qo�r_x��Ɂt�p�?�2��,��(0�u��q8���#QT�O#�Ж������U)�y1J䶲���xvF4�棠 *�@
���pa{�}mm�^��d
�.�.�z*q��D�;8=�Ȅ��*�J�;�8�5Q�>��*�1� ��埻Ǩ��c�_k����L5��hbE�B�����3.i��b��h�7!�u�	�&W8"{502x�؊��t6��U�/P���'63=1K���4��B�l��#���vI�kY�4����հ]|0H�}V�u^籇��x))?%-t����6���\�IJ��Ls��P�`�h?��C0��n�`9�Ȑz��y�P��!�S�	�@t��<6 �VH�?�nJ��i^��ҢX%]��r�p'XBvz�㔍�f/|덬p���M�!�ϰJ"32���� �g��(�_Z��]�4�7�?:.��V�AS �y�����Y����8U� t���<��@PX�Zo
V�����p��I����g)��,
;(�M���l��<舺n�ٜ�[Z�4m�垕����SQ���\#͈�����M���V���O���ZkŃ-��T{�cs/7�1W#�{�v���>�ڏ�Qj%�O|>ѿ.�6a�=x?�`N�Dv���c�c" I������&e�J��_���5�12�����H%��a�� ��z��QDT�B�a�J�=�(���������ZXp���'ڀ�`vRo~	�_%y �Ud�n\�4>5R�&X$C�n��Q��Јǫ�PG����9��Z��U8-ȑ����K�t�񋋷p�aL������6�*��ƽo߾e,�<�~� "��y��J9_�����%�uۧ�$�3u�<l�ε�P���Ye9��;h�7 A̙�
�h�oc��������A����,nc�`�!�(��T{ش�����/��cF[<P���3���Ʈq⚂�K>~V�JOC�:R�ƪ��PDb1I �;?[=���*����
~�o�E S�Y������l2���z���/ݾ�^Ͽ'�r4�~6X��v-��o��}z�����ü��p=K�� �	��tk�1ɼ�x� `��W�}"17_O�����L>�GH����%�p~xT�q)��\!ۧӛv��V^�W��ɉ{�Χ��o���V�h�%9H��ѝ��!�)il^�}������yd9����n��Z�o`����V�j�˿J�C�M���Ǥi6�"Q	��'��0h�	]�>O����H�&q&J/��j���*��i޾zI'�� ��w����"��}�[E�V]���7Uk�T;���-2��e㴏�r�űr�����fa���t�D�v7�F�tt�4�D����쐙Z+�s��U�[���[̳~�|��D�(!t���CJ���5���x���L��+
�Y�nE�	���au�$�fHH4��_%�d�UO.^���lls+���Aꎯ^��.��~R����<�iԮx�P�IZ���Q�R���oa܍m��������K�b�k�D�LmrPμ�T��>��a9�g8 \@�s�K��ٙ�x�U_�i5�#�|}	�HRa_���øv�sFC� ���1[���W�}��=�rΉ�*��� �dl��X�`z1Dc�>���Q��a*lia�P��W9�|��5^�n��+�ON�:����MJ��*���X�*�"�w�m�'[�;`�֫�8q,�c����&�f���;N�j��<l�4�w|1�oz����/�}xd���hA��$W�\�F#��}t?�.�Y��b���b���&[�t%�8p��u�]����w4Z���)���l6� D�,ծ�VP'��'?h����X���b:qɩ�A�D���F̼ؗ���DD
��q9����&U���K�i��vӋ6��� �����=���������3щx9���Z�w;�Ѓ<��=���nY������uĔ���>_��sq��c���S�����j��Ϲ|O�^jl����'�&9�o����fe�H���d��ʠ���q�D��L��n��"N�����6��DQ_ȌL7�N]��g���k�r���+@���{��殳�b���~���������^��엌\�Qo�"�Y.�#M�L�$�?[{^,г��kM�q3���t#��k��C�ӿ5~BO�A��4�!����9�d+��z���V���e;%�����6�S��V�]VbbtΖ^��΍�������[��o5� �6�=�G�^Ҫs��k�e~{��[�X��h~��r�g��:	ۍwۍ��o��;F��Ң(%���sk�{����g���K�05Q�w�b�8|��t�����-5�c�S���{��?\��
��;�P��;�L,�N������>O8����Iuc�^{RL������������Q};���,�ͻl�!N�ܰ�׃��#|ʧ�ӝnt�O�tX�,>��a�K�&D�Fn*
KKCΔ����!��z���d�,D�	�L�`���6��Xk��;2Bl2-/]���"k��lr���VjV��ږ?�º��4IZ�'d�L���β������{�eJK��]�l�ů���s �I-n��������Z���]���"
�d�(���Lj,����b�A�Iɠ��!��u�'	�L�����#.�����������!�6��Zd��m�w��|�ٽ|j�7��UY�4�m0"�򃃽>�bd��]��n�ڷt����23(1`ⷎ� ����^%�e�p}Pݷ<��Cσ���
N�j �_wyu���;�b���<F:��8��2�����牓D��	O�^�����nx�s��˥��Ey��.N��6���o�a!FI�e���q�1HH���*���3/�{���,�ˌ��Ѳ�q�\|�T�5z���ɘx#�i�l΀�Go��/��E�[�*���E�-1��-�tE˿�9I�e?v����t�jT���/#mҨT�R�a�����[�+
�հT�>������bQGEC6�n���PGn^�I����7E�.�S��k�],��{�����nV"�O�W�@ YM���∡6Ĳ	jdes�Yo���8��ȨC�cE=|G�l��ixe]y�7ˆ5������*���B .\Ʉ�����9����RwX2%0	'n���G�?��K���y��Z�$�1�s�/޳�
#觔a7�8�D��!�P�/ѵ����aI"!k7�18�x��~> ���j����`�P�����%u�N����`n�O��?vC9v��Lŵ���9�4�^D:��l圼�pj���q)W�l��D�2jmfE1T��ۋ�@��Ţ?� y��wL�_��_�����b�,��G�c��[/^�苤�GM;ejf������@�s�[�L �����h^x�?�T��`v��q5`��f�&����r��:Xp��e΄�n�?-�Z��]�5\����b,[�Ej���ױ�FI헪_1��ɮ�mlm%�/DtmA:γ�NN��݇����G���-\~kC����+P��~	�����R��4 �כ{%�<�_�����__��ԔD8@��i<�2��������������^���'��GKAl�U��m�Vy`:F�n{�B�]ts8~:�[��P�^�����1<�jJ�rҜ.c��,�)Hi� |O �6���ݥ��qNZ��z�
�������N>�c8�g�?[�5jSl~j��I*�������s\nk������س�#��)����'�����E�5���'��Y�0���4YYcG������c,
�}�d[�񡟔����J�~ۡ�w��Ң;"����D=��A����xU�q�ř�o5әW��E�:�@٬Z��\p�R!\�����%H&�v��.#Fs�J�:M0Z�ެ���.�����G)�dU�b��AD2�:f��9m��4��o����T�!H=4�6sm� A���e�eQ�I�sd�y�F��"sa�ދV�\t�A��\MY$ʓ��a��(?k)��m���Ф��7����~�)�ߔ,����z$��[��L�Z*�>�ǖ+�ǣi�&����$**�8\�O�$uۆ�rg5|P�ٙb��avF*��V�𾷤����[��P������`�Ы�$����&�s��b��S�����Mxg�1*>�KB�y}.�ȉ.���e:n�hy���&�/�\�(&v}��B�j係��L��Y��wɖ����w�f��o-�
��݋��xlұ�iU��Br��9|����P��[���&��ϵ%{�a��1���5��9�_�,�n;�jA��LOr�O�d�x�y����w�fҵ��V/P�>�xתJ�m}©(�?���Õ�҆�{`N���z��_/�B����Q�r{�K¿K+r`|v1�xv<zi���0�Tv��)d������a���Ǻ�NZ<���c4S��b��'♌2������;s�$�OM�ǖ1=kv
���g[9���q�RR�
CϗM|�v0��K��i%]�^�]���(�nf�B���A�q�K�L[]8��3Q����l �cы&�_�J�}ٟ;��\Q��@f�OZ����ĵ�U�ƇE���ʎ�t��f��j�:݄�v,z0��(8Q���l��{<�(;��3��7��ٍ/!�|����Ds��S��S������Z������C�j0m�r�f�a���h�d5RP� bv)`�|����U8wlV����nˌaK�Z��J<�K�\���W�jx�p���t������3��X��d7�y��gDS�G'�Ⱦ�m��7;;.�q߳�[���X�)z7�������`��r�"9�C����%	^�ꤞ�t'0�q�4坾���9n��i�Ւ�}h�#퓉'ݜZv����R���Y��-��4�z{%Y�g=���C�¥�"�͓�U�
M��/����GH� ;MH�:b�y�[�rH�к?�#O��A�	xgJ�NǙ61S����a��4ei��I�>�?J\��w�
�3�f,�V��W1���@���,%����t0����'���{�O�U��!��-�9A���}Q�p���U��P�Ѓ^K��bR���z=@!��1��@�	���i_�h��$��Ԣ����pɪ~�@�����f!�:N�@J7�N��������- ���i����O��.|5��@6́�o5��A��P�7dIW�E�^(�jқWe�'�ņ2�R�-g'q9�ECGǺ��,�8IL��t����g��{�ˏ��VS���h����=+�m�׸��,���i-(䀦{��򧒭����v�;C�er���[Â��2�����ى�O+�U�^{}"�!3?lII�b%*[Y7s���#����<_C6?K������`&+��g�;�����Q��ok<Xl�Pl�0y3�\[����J"���Ն)���݅ub�	k�+�袲�������X'����`J�u���)���P !��Qt=�]Q(���EzA�E#)	���@C���;|�_T\4z�,��Ƕ�0��!���A4�l�0����q�6�M+~*����"���П{>��Fo�Ϝ^�lw݁�n�ġ����{�ܨv�&W��r�l��vj܁�����sG�4:,��R��Z6
��o��`�� Q�$�Qċ�l��A�u�4!^�/7Ӏ��5�&}�I	t�G�>�k��&��{2[���g��%�y���,{b����b����mF�I9���,��Ұ�-��hf�D�\���b�����ƹ��5��gq���t�w_���`�o���z4	�
��jЙc��W��^	��
Ac진�[�֏�CD70����_�-wA�7����W<����g2Ю�Rff��{����4H�DE��>gK�[ނ&si��1��X8��~]k{�hh8��n/��`��,��{�[	�^p"��~� �ށ�v�VC���"�u�{���G�;�m�t}D׌s,Ow*˽K���L)�|�G�_K�	��i\����r��ޣ��|�~���N���ǩ���K�5�f�p����qh�,��e��gv>��m��8�'GGGW5�� 9��\�7��7�dj��L;)oOݻ~�Qh ��������y~.o:�N0����r���z�/��hi��3lT�V@��}����(����8�U�u�����Ӗ�ֿ>y�@ڤ:���,��yWD�@��Vx���/�R����{�L�a��i�n�>��,� �@����*X���eT �ɨ��l���5$����0��8�e�<D>�/���4^f}��a���^3UD�ǐ����	��Y5W�];�E�Qz���HWEg������V�;����C��'|�[QB���� �e���f�_*l�:}|��>`�8a��w�
��a3�
��Y��0�C�<���W����0�;: Wu�d�Ŕ`�$��SLÑ ����C{��$�IG&�M�̂�
��������4J^��&*:�FB'RRMG1 l\���5Ϝ���R�n�����K����5��ӍYM����z����k��c�lѿ�����7E�� �egc�������2"Cq�7l��D�8�B�uW�i�|)���[
=��J}h�����Vsy���J��khzz�{�|^O��ʊ�atola�Ic�����K��-���\��o�!XE��8��<Bc�_�(!�<ԋa�����������P�Ƥ��Ԅj�p�]|x�|���{�:1SE���TK[�������f����~�����?�UJ�0�hGݚt�����N�a]�Ng���UY��`����?�3��50�0�P�.O��8LCX����%ټ���Zy����� �4J�_�h����#��[�H{5��������Y�>��k��Bk����%�^�,���2ؽ���m���2E��B���UGR:B$~^ �� Z�^�ȑO�V�k̯ǡ���r�%�<Z����p\l?�Tl)�<����.��� *��!�;��U�I��lo!-Ymq���YjR}he�����l+v�@a���o�5��,��.�Xg��M�ܵ��^���I~��[ _4�y���o�f�׈ȐH>e4�*����/�Ҝ������^K�h��{�>䏛⤊�*I�UP�σ�-���,�.z�6���3fh��ڠO�ަH�4;��y�9R�Z�����C��t��iQb(gf!(�1-��4��s�G�N`�� >���_���)���7ǹ���9M�o�����U(�P�wA��V�[��PP�F��Y�L!�5��Ld̖c����!��7�=�f��a:^�}O�����T"���%���h�'�����G�s���M��(,I,���I���@op_N���c��-)��8���\�36^�%���w�a��ш��v@���kK��7��2GЫ�4p��\n���򭭧�ON�D&P�K<�d�(�+DL|P%e"å5����LnE~���Vs�ģHH[� }"��3_�n��?y�E���f�֝�oܕT�.TsX��e@��2s�3���wZ>��s���-�f���U�&C�
_ΞT����Hc������{)&�:cH���:esq�ۥ2F�<��"�>Xa�;�hQ�P�8P�4�1���'�W�Z�*�g�xE��M�w|��c��g����0s�\<� 1�?D�Lcs�D�x��9���S��.�<Ċ�g!���Y~�G�|/�uX��8ؑ�����kF0{��祪o��u���.�J-*M�v�MM�p�S��R�no��&�Ԓ��S�!9Ck��y�-M���bH�Fr�ڝ�P�a�׶U5a�z��q��0�.a�w`���ܻ����A���І�d+p�M��`���o�C5�k��	��)�6�XѠ��8�L��]��Tv�o(|z1�z��p���9⍆5�*A"ey��O, ��Q�?4�0�oh2L����&e��u��'������R��G+���J_A�Fצ�E��.��󦾓a��F)�|��`r�%�����6`���]}3�^��f6;N(1�ְ2ZE`*�pA����6~�R��pϘ��|}�h� ���d�Y}����F��֋��*B��+Blfz4�a-ي
r�^%�{sM���^J��F�a�U�����[҄��̀�yإP���Uآ�jj��pn��@2��9����q!��o�l<�;n?u�̏Wc�j@�
Qw�;�#:�j����r�_����/��������rW�A�,X���gC�R ��1�����UeU;�}үa�>>4����q�6Ta��� I����W7����8�V^(�(v�=�WIup���$�Y�3�b"�N@t���}���u�ͨŜ*�#p	y�"s�-m<|���yy2,�'�M<�L��,�F.÷l<j\®6,i9]#s)Օ(��(�.$�P��� ��l\�ƥ>�����w���"�xH)�MWp�c�-��^����M���C��77�h�
*,x�Lz�(�N��dG7G�/h@��GXW�?��,�o$�b���I0V�T@��[043�f���w3��_)l:��g�_iU�
ϫ�U�w���X�	r�@X��RqC㫔l2�|����k$㽺����dl��Cc�i�~�p���jN�*N��Ď_����k8�s�������@a�L�L�.�7��鑘Gi(>��N�gE�0lu�x-�.:�G�ò!,
��Ñ�Ru2��fl�n�qS		]�kq�s���)�Gs��(�Ix�d�B׺������ w���������t�=�Tܸ�f����ݑ�C�\$v'U�Z�OԕQy	A���B|0�9G�9�͒XN6���/��;���?�8x֟u��r-;p�dd`[?
{"W�F:M�jz��a�l �M�(A����b�݋"0��q��`���
�-~�Y⡣�1�/������zXz:T<ؓ�S����;^:�߱�v^+��eLg���H�P��5ֲ�4���=�ki��?�z����9j�·���nA�<=i��
�Z�(���7>7K{�H�sM��EQ,ݪ3��ЭtW-z���'0�F:����8��6�6�Љ�u� ��4}� ��N�{����,,C"�"�� R⫎�����D�Kώ��Y^��WR��^T�Z�?,f{��0�pq0�1��vͭ�jt�~ڝ� ���
�0�^��Ȋ���X�x`��$j���1��Nfy��3�g�رz�듆U��=��E�"��v�n[^h�j[f�d�]�h�̑��)�UVW�}�b�m�I:�e��J��B�x�1��7MWt\��4���-��D�ca�c��u��E�{�.�+�K@���"�� ��Z��xV�]���̘���w>g�f�[���[�_��F�Gm��?^P���x0:��N߂��*x<�4nh�Bw�m�[�1�Y����C4.�Q��}�H����'K�7�+"�8�r��W	X���#�œ�Y���=ɛ�4W�
(Kf�)��+�E�񵂣���{��!���x-��}��~�d+W������<;��n�uR3x1��VTt�Y�J��������_x��ɏ�N��ة:�I7���T���v��f��7�y"SrR���̚Xt������vKa����K6����eK1ob��<�F,+�k:��l�q=|J��l�bi�\~ѯ��!�ى�HsO�w��M�]�)iB���";Ylq~��r8�G�p*����<S��� �tGx�20�0�S�Sy��G����>*��%��pf ���{��j?�)��: �ly�(�D�=R�A��/Z;�EgQ�[�]bv��|נ�u�?�"�ǽN�#��={H9�������ǰ�$}��U�V4�]5ˢ_�'S���q�L�����c�֯���Փ��X�ɭL��U���J�3���uj*�k�����lk���n�z��*��q�l�l�E� =Z�ڤ�_�j���g�)WR�q�����2d>�o���K,��ތ"�K���SpE�(��ޅ�dHN�,^��5�B��0ē�.�����+"�9|yk8r�q�]�Lנg<�/��b������@ɀryM���=�Z��7�p�+���Y��Ր�@�o��2�N��=��nf͊xq��7�lF��`ZƆ�(�����2āi�!ƫ��A��p��
�X?�e�X�����D��%s��~�ƇXg{,���	��y��zk��|�w&�~e��[ ��ձ8�C�7��R)/��\�)���*��GҰ5�T�����St�^�Zhd&�͇$񫯢�/��.��ߴx��W.��d #IҊ���7�������X��ֻ�v)a�E�sih;�A<�3�U���빡�NI��$n^��V��¨@Rb��sK��� ��\E'ם��UL��L���O���;���6�I ������{Fx�Cȷ57h�a8����{�C��Fl�	O�.`G1Zz��oE9"�v�si�m@����O(��a��d.t��A��1�E��w/�3$�G���@�k}��"�ieH+5֙��
a��=ؠ�oX�R)�����5D�y�3{������#���e�*��$����a7�/�k��k��C.cƸҥ%
v��N�^����鵴w��_���S\V��]#R��	4����Ѥ0�p�\؇�ߐ�0u�e�m0��qy�pO�Dv_�l��YWކ`��ӽ����۷5����$<����q04P���N�d�v��{��v���0�~!y5�1���Q$�U�V�"�X8{'cT�1�d� �zu@��Wtk�O������bo_	BE������p{��_:~= `�hJ��a���]�'�ĝ�������d?n��T̖�·
=��|ڔo\ۨ�"�J����w�wv�*FKP���C��3[�2�(��?�_�,��R�T�\�^}T�p؍��\�4)Xr=Пu�BF��UDM���)�z��mj�n��� ɐ�V�5�"N���\��ֲ{���r6���v���l��K��vя* �}h�4u��/b�m��W*0��,��mvB�.�VZ�E`�4�Jd�S(eXɖ^�o�R�O������
��l`r=V��Tp���y (٧���.{Q�^U�N����b��z�W���t��E��>p)v��<`���4�3��vd�W�5l�b���:t,�J�Mw�L�H�Pg��Y�r�{�7R"_�δ����4�~UBӼ��#b%
���u �����1k���9�в*V5G�[�C���9�L�\Z�g3ϐ��ď����GS��pϻ�N�D��L���GQ�I��>X�BcU�o�:`�s��"p<,�r�|�Α��@>+�i�I�;�����R��.���q/ڊX��RΘ��ם�x
+/�\N�q0#�OE�{Od����h]b݄�f���{>q��H'��!�=�Em�}������%˙�U�̠�G?!	(���a����)�u��ڮ��p穥ōp7&�Q/�Jøz��!wTl�;�x\P���ף3��&ܙ��ƵOz����A��ӛ�Ze
bJҸ�*���s����xˀ����;!wiq���P��E�CqB��-^(^���Iq�w��
��s��}�{�aɗ=�֬�w͚���Ʒ����#"?�i�hHݢ��R_��9.�bؿ�\I�7������yb�<��<��h��뼍p��	�aS����n���y`����q�(I�_\C����[�(IZ�J-,f¿��Kܵ8d[��2��mo��ʽ[m&��|5�1]�����}�O��Y���i+ A"Q[^�E5�yl����RȐ]V�7� �A9�fn�%e�z痞�Y��h0B���EĆ�t����� ����A�_3_w2���+�S�L���te"+�����rl��]��bj/�i�c~���B��5
�j�m�!y0�lA�z&~�����'}�8O�^8wk/�s���	��f|�Q�xw��s&8T/��j��x���~\���q��ܑn�X���\�C�{��;��%��m��)��D��$O�N�C��/����xFˠ+��ǆ�{;�܇�̞�����b3[�u�߯hh��b�+j7��ޔ�~0ꯏL9&���҃W�z�|��Q��i�z-V��6����؂uST���?r��n�u�`�uvη��=���p�i��	�}����~o�+���	.&{gGV}���o��ơA����P�<���#E�9Ė�^�(b����W����ɲh��C^�?|{����q0��e�>������������ې��S휚��C9krJv���HY���X������X��g4��>)�I��>;�߿���Q���t�v7���7��!��&vɞɀ�>��M�����������N"������2�\�V�M�pY��ɑ�<==N���u당N�]��*%C�j4�CBFRX�d��-�=�K�U�-g�e�vr@XTt�I���f��aĦ�Խ»��%���`���&cU�e�j���sr4�)��~ oØݏL2�t����l�LI&��j 6c�+$�avc!���%�C��cw��τq��q!RkJ?�V�!��yԞ��$�`��W=ܽ=��
�^�4Oy�
/n��7�[k)��԰�̼��Kqq�}֑�8֗'UfeV?l�x��J3��?C���Ac�<��6������7���!	|'�']��uV�����t�2g��溁�f,�ոH�����>��}�s��lL�ꓲ6�]��B���-��L�����ad� ��z\vj�K� ;Sg��@�9/2W ���]I���{��56�
G���� Ά�!x�y~����ք���~m:��%W��O��3;�,�ʽ�U{N5��z>W�g��j��;�wf	��?z�"A��6������#��SDN�D�ø���z��nάq�݇�/L��i�At
�b5�U~����a�,?�ⷻ��-$�#>��f��8�Bu��y�I��"�����v[uEC��&�u;]i���#!���8�[|X/�NOx���_�պ��jئ�2�2�a�&Ӌi���bO��#�e��#�ҫ��!�,2{OR�B[���V� r�ي��IϖwU�@zs.�I�C1��" ��c�%�:!O�`&�I�����q!
�`05M"�"��/���Khw^Ph����MoS��$��(�%$z�4�$���_�z��필�b��v8,Rw����NS�I\�<+?LÄ�@{�����x3]�|V��`�0_bV���'��
�}36@*fd��c��`F��;|E�T����H��|;����i@�1I ���*�g\ɢ�'v��xY���V 
M��`��S A�U����w�9|�$ru1��/��j�ޝ&��M�|�	
Jѽ1�ӷ�᜿ M<���Ny�a�"�b_)���y���G��GSI�ZΎpa��/�Ȱ�>��r�z��.U�<����$�� �cX�>����f����1� ŷ��;4_V~���z�z��	���{�󩙌 ��j5�L�e�u�lS#1�X5�
��/d�ih�$�k�Ze7��?�BlWt�Mߺ��"8�'3k~��-����vu���{�n�}�s�9E�V�h�'4h�rw^89:Rg�=��ؐs
1���6z�T[���pX���o��lݞOEtA��j���HS��-5o�	琟t�*�*Fu�Ot��kr2�����cL��t���Ս��7�g~@�҉�Z����"���n�"�B�k�MoD�r�R��I�O/~��X>�V�"ۘ��'�����#��'�)O8Q�W^��!�h��CO�G�����J.��i��߂��T��g�n��&[����x8~�Wg��� �>�D�H�A�_�UJ��Um.&��g�� Tl@���wU*��G������̌��[ZG~cn�/��bt4���q#�*E,*�Z�g'3��������D����~a����Q�Y�8w��Ӱ����m,x�/��d�k�RV���@d��q� �����;�$�,���#��@Bg�s���S%x�T->�7c\���ИZk�J��ί�h̤�Ov��}8HDS=�3�l�I�q6}�uz{������t�3�F�Џ��<=NvD��:��ٹ��Z{��5)��ZE�>�w؉Ǚ�+2�S\ct��
D�(�j��l�YD#�����okD?r	��E���	��&2��ՁW��oV�mz��~ŧ�b�G����@�)=9�4Kh��	�����|���:{\�$;�M��V�{�#ҿ�x�g]�K��z���vFK�),|�0�1W���;?�v3��ֵkև>����/�o1�j�c�4�#۟�(VclG%܆ۂ��3�Ê��L?C|j��c�h$�A� 
ǲ�8���ϫ:�t� ��x�1�h켺�`@��Y�T ��u}��+^����&޻��ݗ/j'b��p�M��55mM{� vv`�.LFtRz��&��wj�c�x^v����W��}(�N$����Z>�>�pK1J|n�=C����W��H_c� H/�޽?�9�ڛgxk�QXY��D'p��Y�.`���mp+]���I1�IY5�49�|
b�߿퇽c
��Ri�����c� ��eDI�5Iqz>j�`/ݵ��c�6o��7���O����x7�v��_ ��c�(蟯u�~4�!�=�Ә�!��@�r��Y0�E@M@�w�٤{�����i�Sq[�%3R�{	�ޣ�w��H'U2>��䜃�t��7��J(�E�=ݍP'U��K�}��/{Y��ޑeA����|6\L�y�r�8^�'}R�V�<�n,�uY� �ȭ��a�S֦�^��|����ס �Y*���E9:�޶
3�#)W�r�N�Tť�;W�Ӱ�Ƞ,��XPe�9V���xqS�nD=%��%�?1�m�e��u�n��?6����K��7�<�i?j��%)C�����Q�2����W�;���|7,$Q����˕�-�Z��D��9�6�[���e�m<�z4�SQ,4�5V�vy���d�"͵?$��a�ġ�L[E�(�,R�������[�c5�U;�� �#��ry��
;�gm�@N��I){D���'z�Mo��������o�(Bb�yb��R�^#���L�nE����)�Ul��Mu�u�h"C�ix����y��n�᧿;U;XX��LL��d�,��N#�fQn&|	AY�#U���� �'M�O�Ϳ�z��%�a�bBM)�o��t�-~X�_mf�+J��A�q<��� �c��c��z�4
�e3���G�T�yC1I�X��ԧk�ś���cz�k�HI��k
F��lHm�-�=y�;)�O�)����
]�A��M�3�7���N��zz�UTͧ��
�/d�:��U�~4�%E���	.w*
KM��wb��k�B�</Z3$1ŗ��~w�Q<���NPzȑJ���f��qQ�2�z��=M����۳�?�a?�c,A}{�6l��Q�?g �-�|��v�/n<��3�8�)�"y������@D�pZ��N��b����q�_MOޥ��#	P��5����WU08XJI!ykT�/�q��{������ك_�Uˑܝ�� �YИB벙����F���Qڑ�O-k���BX��79����Jʊ�e�γ,�\�� iUG�@쇯�YT�	w��Q������O_p)ڦ����"I���ƾ��lN���k�HR�吋�v��+�ʹ��Hʉ�k�:�JQ2�~�|��:x+6�lo_�:������J��@��&��G"�n�'��u��ȋ�GE��V��x�z�bY$^T�1?��~SsF����~�=F*&� 
ls�Q����>��g�p�s~D��ʃb����Pv7�g̿gS9I�ї���Bς�0�L��F���?���E�I�'�iZ_
(����������eW\ �w+Կ�F�7��;����N~��0����E�������΂�ˆ W' N�a�V�Å܅�k��G�k��a��ݒ���§ʠ���ҟv�F?��ߢ�<�r̿�!۟����'f�4�[�����w��:=����b|��2ڀҔx|��Uh��l�Þ���=_("J����;�����������F��п^ �i&n�z���s��E=ʘ}�^�f�m��lg"u�J�w��H��q�Y��}6��eE!d���xjFg�`ֹ������#E�5��ð�Zq}dJ%�:�x�.)�
��m���L���Ǧ����zv����$%d���Oj��ϫ>�:=/V��OW��̡�,�L��*����wH��{����vn�dP�V��\�W1c(y$ZR�F,�[�#0O�M�����
)k�yqñ��?ô�:w:�:��R�i��� ��1�};��L���������ʵ�⥲�Y8�g/���4*~�G����4�Ύ8V%kʘZ=kU[M2\�GP�B�u�*�����F�F��G�?��h�P{Z�c�[/�D�����CG�I8�47���I6[��|b��H��BAU�)d�q�6FZ%�L@��M�萋��{.m�~�N�>��z5NHH�a��	D���C.¥͒�W?�vq���ɄU�u���y���H�[.#�5z�ݟ��xfD̷�Ae9�a�?���v8����*�EP�]"����yK��U��)j�� � �$ �$:{ ��X$�]/�5C�>��J�vq��B<�+�?���̞��Vn</ax,�{_�.�<���W��Jb�܀�ޣ98#D4Jf�`�L���H���5�T��/ڭ`�2�*8<HB�R���b��;<)i���	�7\>�^�Þ�{�����6�5f�<��'�u���W��Z���=��ȼ���b�)�i�0���!�Hd�>B��8Q:xJ��B�`�`_�؉u9��f���wF.�p�?��O*�#��4Z���}`U�{_k_z�0Y4"����Qc��䐨���O8���=�y9��I�6����fօ�^(I��4G��F�T�{|�¯*m��k��v���p�h+W:�)�唀��Љ�u.m���K�͜;E�[�Z��*&��g1>^
��Ey��RF���䨒C����%�>n�oQ8��,[��l<�I��bɎ����oX�v=���T�p��Y���.�4M�P e1ׄ��@X���Z��/��ө�����"z����K2%����ki�#�ZI<���:D�-/�g������H��b���a-�S��p����&��9�A>�sNiEEw����t�s�k
-�����-�P\\�U�l�?[��M����oڍ�йR(o�{폗�9�:�L|�&is���N;q�n�z�ţ�EA��I�P�.N"M}���u���B̶r�}5�RtUD�^�f����a��0��0�'�������4{�=�g�9M �!X�X��A�x��r�}��V�*ԕ�%䑖��=LB��������WZ��ȕ�lo��5��#�ـ��[�JSF;����jԉPAE�o����q��u�]>�EL�����޷䬿�𛀯/�MM�w��Ƥz��L"�1�="}Z���Q?�	ռ�v�m�9v{o����Y�c�+tC�������q��c/.~=Iv���R
�ګ p��P��6$h�T!����*�Ѵxvk�jN��8N��}>��=�B������f�t�Q�\��=�N`�zDX���/�}�Q�T�.�)�_�7,�$�_�f��Y-PBt��A�ߟ\ǩ�Y��Q':#%#�[���jmɼP��<~�������o�/�׽k��/�+�}5�������}�2�;�!��@�o�**C<?E��U�I�x��
�
��M��ssd=}r?+�H���tB�o�-�;@s͟Y�{.�Ϋ�֭M�4������<�N\T�u���g��4:o�w+���Q��fi��=?���]ќ�S�_��e�$d>#T92P$���ȿ�9ҍ�ir_;�Z�)���ְq�!}��pn9X�'ȼ��4��U޼|��!-��w�z�������c�D���ĵ�<�:ÿ���uv=Z�}>��?�u��)Ǣ��	�"I$�)x�����wi /.�i�Hz� �Ȓ�v��*��P�n��+j����y����2Օ���D��~+��7ᤊ�ު���fx�Z)F����ʧK��<�����k4���g�'���8�>
�	��Jڦ��D���n��x�B�θ�)bXʩ�d�=�Y����v����`�-A� 8�)���(z9W`̩Z��~�l@�"KD��ɥ��	n`�3ka�em�$���\L��~l��(y8��r���f����l����C�J�n��Lt�)iW_m2�<����24'gj?�C���)��l���+w�����^��ޛ��w�/�x|C]	�.}Zt>����!��|�����M�}����$��ßtvy�f�편|���5��s; �����6�V�������N�y��ڧ�Ō�hK��)�n���+���y�E�o*K1_Jp�����<�������h9vK6V�~��/Y�͕u#�Gr�g�͔W^�D{9���3�SF!VS,�w�_?h%(�X ��� 3W�Q��;'+|)��J{u�����o�\��!Y�����n�դ��eד]� d��� |���=2�4%��=�Ռ�K�P�/߽t��D�E��p�R�I��jdK�_�>��i�Kf�n-�s/�[�|:���.��vO*���0�܌]�����)���@c��U�Օ}����CbU? ���W:
�&�x�g��?V`��­i$����#ϱ����s;
<3�8��pwi��{Q@�v�0�ꮌy�QG���C����C�"������Yۊ9��"u
�3ф����д���(釖���L��?����_%E���|B�a��R��t^���r�s>�h�sD���Ai��5����i���"@*�B�C�1�p��j�b�W"��23;k֟E굱l�Q�#��|[{:S��-% 6e�P�G =|�ڑ��&�tlϥ�6�1����fm~�����2��N6фʅ-�`Ր7]ޖCm�~E7BL�j!O������Tk��e`��
��;L��,�Cۂ7�[N�˺˟��*_ɠîs����)��k����ζ�)����
�(^μ�*�V�ZB@�x��Te�AF�Е��7|���U��o:,��Xؾ��#Q�����]���)>U�t�׎����V�������e��uƠ�� #t�8�wOߕ�F2�n9����?�:?���9�"��|�&�=.�P$�/����!�S	F�,��i��X���NG�:��AF�(g}���tM�{<l�s�m��U�XeS1�
����}��wH�=�Ʋ�%K�OY��߶[��f��O��p��x_�
�$�����:��cs�LLx]P}�� �#/~�C6���)!��p�r�)=܂�2��c�l�:{��	KZ�J�t���X;����~��K����x�G&ɇ�gTbf��7�#��H8�G��o.(���ey"��y>$]�o�i?�#��U�����n���� ��>�#4$��T~'�dWxC�W�s���;On.f��S4_�����j��[u��sԡ���
�Kv~�Ngr�����Vk�Eu�>ڿ=�
����#��)����1����F^���7ABp���^��V�?�Ѕ,��3���Ob R����M��F4
Z#/w��vj4�Ee�_���<���I�ZG���z8FX����#3_��,R��\1BoU�v(�[+]z�
���$�~��Xs���U^�@��5�VL;K#�;J��@7Z�5�<p����K�4���M���彠�X5�8���#�������*}��uУ�cjI����~�����-m�N�n����{&�Q7e��^��09<�A8��q�0���3B�O��Rr~��&z7믎�	�=T^%�U������j�.���.��??��c��#h����H�wk�?���#����lx�.�q2�( ����<2���9e}��>�#@e�JR0�K�3��;5�ùP�uJED�أVM��-Ǉ��'��F�(DTޫ5ͮՋ��N3������W�\p��M�a)9�Ab0'��^f^(&�S ����>�\�P7T�0���`��jr�jO�d�̔���z�N�o����zO���L�,P��{��A������jqI(�����
����~�T�E�0-�dI����F-�BɎgƷ����E0����6�I�w���S�`��?כړ�..ђ�����W,_�*�7�T'�c51g�9w�@r�O��7=��ܯ�=D�u'����w���/k&Ó�H��~�2[�⶗����&Z恹{�j[�����~�������N�q�\��CE�����pO������]�	Wi�;GA�.B�^ID?��kգ _O@*���V�!���Q�q�^H��S���P剻��p���{}��dx�2��^G��N�~I�P�V���x�8�Y������eHͷ+5`��\�QP��뿫G"����3����6^�g:l8�L1fB�ƽux�x�
���0r�-��<�K ��PΑǖROMM?J���wzf�]>�<���yM^	��`bYk+F�w�b]�l�k/��c&�ر�I0r���JO3��X����?��'��5m
����p�`��))�v�$q�7�-�_�SG�^�Fr�؏}g�w��|T)���� 8�Sm�q8�>z��K�|6fG�C!ފFJ��+Hԧ���ʇ��.�������8���<����\����SSQ95������.����S���)Ȝ8Y��Aٵ�༿�G:��.M�n���\]֓���K��c��KL��]���sQ0E2�{U��h4췌j�1S�b=��{�R�cw�s���<jq�P��X�y�dj�w�Y�|��{>�����^��S�����v}:�l�:@�#�WТ�ִ#�4�a@=g���ֹ��qȝ�����q�E���jL��|��V6fZ��x���"e����~.�7���n7��>Y����1���W� oÚU�)���J�(u���e�G�ϼz��in���K0iߤu�WU���}��?9�7�T��g����e�zVyOve״�����U	m�G�I�q�1�x8��^��úWQ?�<̌�e�D�gdj=��*���f+Ycrm��7�)YǄ�����'z����N2�ZO+�$z�g�3W���h�C�j�B����8��rc�J�mf-��'�E����8�.���B̿Q.8���3�$QN�恽��DO�8S���&=�B,���Z� "�x��������,c�ǒ�I^��i���~�lؼ��ΑQ��*��L��D�/�j�Z�}F�4��T�h��ǐ3o[��pMN(2�G/�&�d�"�x�ј���n����Bc�%>5���/\�@'J����LV|�Ϳ�+��u��j���'O���5�!���/���-�ȶ3�j!�w��Z�d���� ���X�`x��Y��w���%�Z}�k"��4�6J;�Tٗ�1�?�?�5����5�`�@��\�FV�8]͋^SArE�ц�h��*�t��(O�	B@Ic�>�1�E�F�������0��i�S*����[� z')��	�F���������JR������G���ג�^@O5�G�h�G!���öF~��ߊ>�Bh�><x���ׂ�8z������M��&s/3�>��gn���B���Fc�h�I�ٓCX�x���7�S�5������︓�ȸj�Y���^�Q�g@O�O��D�7RǍi�4}O�=���	�d�}�#1�'�`EVUr��a�[sN���`^��?�̓"���j�9+9ޔHyֳn�Y r�.`am^�i�y��%P�Thi�)�:!xɛ*�bAl�0	1��NV�B4YM�jD�ke1�x��O����J����JK{RO
�/��:�֤��}�PM�"�&m�����̵�N��p�T�� ��6�Z��ed9���r�ls�\�7\0�4����_�덩����}J��`I�����8�{���k�"�bd$KZX~O������b3�������|�1>��f�ms诃)�6�-S��O���c4�v�H�Em������L"�@������0˥X�~B���K�1U	C@)TyD�V?����7��e����Y��«�w���Th�`�Ir���X�h���;�?��̒o��������y�)��
�Zq�!vYn9�I�ܬl�wx�Ocb�m����"!چ�QVl4�C��l9��`=�>$��Ǣ�N�`KA�`w*eD��)VA-Adm�C�r��D�:�K��*Ƞ�'�v0�J�~2hp�T���F�H�~~,��(0���CM#cW%�NU{Ei�����	��?�m�C+�ޡ��������Z�Jb������t��S��^��+�W����?gLPL���%n�^��x��>�./.��N�m���DQm����8��0�[y����;�B��N��_}0X�(����&�ʞU�]�N�� f����N��8�əD0�t�D�U�|���!��ɹdO�Z�������:����j��X<[<��q�C�i�i�/�<Kb������b��d�(y-x6n���X!��Oy���%��YL�kD�}���Y��{���/�T&�Pt
�w=;�)�2�F��1:�c7E{����V����=-�O�OZp �|�RLS���R6��ւZ3D�EP*$gb�:������K�	{7X=	ps!;%k�z���i�	�3Yǎ]�0��lWIYds��� 7���KD�t��9�A%���dT��l��w������@�/����l��G���;!�9��q"l��g�����3�wa��/ɂ���QW�н%?h
����F$M��@}��8b7�A�Uh4h�5տ��:�v��f	t��{#�3�^xل���q����!��I�-C�r[i��/kCy�zd�g�<�'Fs�������1�d�h#���.,$��0h��ፊ��%�pN�F�4T�Օ�q�4���[���q�[�g>�x����<pI�?Qj2�C��DB��Q����\����3�ЊX2����x�ߢ(��B�=��u������j�ɜ�P�E'(���	}�.a�Ő�i� .Ji`������� ѽ|�+��P�!��q��ؒ�-d�OgZ���Mbyx�b�;�L���s̜��N�;BR�lI|� �wϖ{�=:]����K��d�m�"շ��X�C
K�UY�d˼r<�^SL�����W�y%(��;o��Wڭq��7ß�"{��i/ҚQG6�\�l�0���nP|�0jx�DS*r�]_8~��]=�"���:b�|�ø�e�6�	!�u2�8��it�K�y)��b�B�`���@<I]���X����ߪ.6�Wm�q���Ѽ{�I~c�5Z�{)�����K	ö��hKwY/cH�3�V��u�N�a~i�<1K��r�C�_������ɕ!f�X�hK����"՘��7w�ǌ]?y�v����(�t�!�gQ�'��Ʊ?9M��f�}��l�wE�mŻ�����S�1�E���Ͷ���r4�9�a��t��lM��o�B�ʮ��K1!% �A;���I��V�-ۄjܚ}[�����2J�ꦠs�~k��-H���	��*��
��	���:m�[����6��J���&���+0���$�n�v|�	���a��[Rcyl�#��T� ��߄oUړ�8k�ڝ�/�+D�9EBa��A������DMb	w���k��v�X �8?��740�(�
Sށ)�(��|�,��s SY�lr���_���伀���҂��@�&i�z�~ylGl���n�s�{�1��l��Y���O>9�"n�C/�P� �&��ܞh=��.ʹ.��~[	��?����^΂=D�&��U[C�5�Mf�����)9���z��O�1$����թyRuhow����J�<�<#gc���?��l�O���&��� N�bW(���fH����W��@�m?��Vڅ������]~'[����-cr!p��~ϖKm?�{|�7��)ߎ�������%���'{����`���G=F�ЗU��aZ�Q���%2��k�[�L��ަ.��|\���8!lp���^�wn.����+O�o���	�Q��� �����>3����޲��Б$)����w6�=��5��(~�䉜>�l�pv��:��[��5+��v�H�eyۺ�r/��;�[�ByO�NT���G�{^�8q�
����톯�g��R�+=�gw���+Η_g��b'�h�v2u�����n�<��B�8�'�X"��kF|;�,���\Zs�3�2�N�j	g���d'L�Bߺr5�c�8��A���ӭ'-���F&�\�%Nio�������J4��k�</�����d����Yk�d�ҹU��ܞy�jˤ}�Rj.�*a�A�V�Pn��	+��f�d�Ԟǒe3<�6�X��.��4Ee�*�qS��	l�4��@ͱ�3E:�y`�1&�:af���;�E��'�-2�+���'R'�����Ҷ���4eF&&�fȟ��	(]N �T���A��2Xs��]�5�ݽ������N�{!
C΄O&f�����s~�1��a����U~4;�+�?D��Q]Pvx7�F35�[�2*�ۚ���v���h,�ȴ�b���B�
���|sVi^�V��zn��	h|>u�ܟy�f��_��ul���͏ߔ],��u+su��S�Fx����}Ez����G�H[71�g�&~7�Ў+�|yޏLn�Q���!2���C�~Q
����!��C��.��šAe�.=�N����R9D޾r��Rr�WX-.�������ԧR���p�1�㠹�����_�8C��-u�~��c5B�#�����.e\Z���ؘ�K���p�K�k_�f^V-�}��A�f���j��N���Ji��IRx��Xp ���	��\L��ڢ���_���L���YM�UAڶ���~�|W\����n�BZV-����S���8	՞�w��~4�P9������H�F����+���%�ˍ431L�
cf�-�/�rPz���(�m��U&�r9���Q�!e�#��c�8�M�Se�B6�z>�~䙷i�����{�TR-|�Bu�O�_E��\����(W�@h��@XN� ��Yٲ�"�.{���D�ԫ�l\��t1�.p�uK����+����p<�ꞿ��n	������v��z���`[�'b�h+�r��S�~o���3?蟤./;��Vtg��A���N�k��Խf��V���2����,�:3 ;�h֌�����Nf��Y r�y�Z��g�;�Zn������I�	ZHuA�t{��|p��KX���,�y7�Z�T��ν��]��LSpo�̛C\��?2��i\�,ҡ�A��.�����Ѭ��)G�4m(��,׶,1H:tq��Vwh���M�s����s�7~��[�S!A=C+������V}wP+x�­H퇒�jfz1V؏d{H^����$�p�Z���ʊ���/�)j�Ǻ@F�.�X@7w�i�L�췖���t4�D�Q�2�-��z��"ʚh�J�9>+�8i�|@n6>��G�4�^?�J��C3t�K�Y�D���[O�wӽtn<�ֻ����n�T+*(:5	`�ʃ<Z���SzA$��<�z����B�6>�ほ<W��:_DB�[9�UZ��/�M��*v���\�|�ѭ������)����^Dp*m�F*�/������04s�������th��^x���P����0"D�"�:O4X91YLЖ)D��D��P���gK��+x7�s7���5l�3��)�cf;���3��Fx���}K�͏5kѭ�x�R��u;��._o�坛!�	����YY$�UB�]71L����]-�FJR�:҂����;]]�OI}�'���\Y�d��Qk��l�&LV�$T�fޏ��J'q�U���L�_�AsK��Q��H�Z7�7 �ش����Z�S�]�G-�#Z^,�N�Z��B��%g�H�
%������U��l��e�Xd�On�E*�KK�WH�S]N�Z7�I�@35Uѯ9����<��|@�����*���WB���,u�ܔR����?R��v�w�KI�xSJ�KX�c��� aۭZ]z�2��S�kږ����ۇf�<�o����Ï����w~"�vη����p~VZ^}Sͼ�
�G��2>�zF)1ށ��ƽe�=��6z&�!��%���󵽄�+�f�޴H6�-W�Ґ��I��ٷ[zd�Y�{)���f�~z0Y�Ӵ;�;߻-�lv����b{0��A	-����3sj��g�-�\����,Sٿ�.���_^�l��ֿ�ŷ�(4����l���>��P������w��K�8�7��"���s�R�l]w�F��4����j��S�O��5˽b�0����Ʊ�. m'j^�q��7{'y;�O�R9�Ju�X�Ȱx[3L߆�4+]ݢP}�"8��c̓��ϝ�y��)���+�TT�jm-�� ���#۱�7g�w����}����;׾6f��:V�=]�='Q�����<)uI~ڒ�-~�JP�����w/]��)�((����<!̶G^����&*�zЗ�ʍh�6n}} �\X[&��"���ؕKt�KT����+CK�����������Q��U�Sƕ��3D�#ƙg�j/�Fk]�D��'467X�8��Fth�W����1Ix��JL�i�٪2�|
��d�bs"��͏ҟ��~�J�v�+�>�r��'����[�O>4��$���_��е��4q��~�\��ݛ�@R_�-޺��T�쩎�;l{�\B?
5!���E(����>S�xϵ2ۑ����k��'u��ų��(_�dgteK�.��2�7e�B�9��W�vf�oW�}�/ZW��(�S8J�_o�>H�������C7���}0~�w�%2*.���|��W¾wf
�P{Q�����ʠ[����٧\�5�TC�$�u��EHo^����4�W�P��盾s7kۖ��`�N�;��}=	8�F��
�|?� (��]��z7�nf	^����wt�/N��XA�|�xoK�doP�ACQs�#�ez@�B��`���,�g��q_m����޻��:Y���9�`ltb�4��g����z��2��x��mh*��U�B���چ~\^�M	�����	!��}6r#��"��6��F$�4ֿ�_;���%���T����c�e�@�|�����@>��˹푀R�[J�4]-~_[�2�v���8��qg�-�qg%6��\Г�1�B����U�ͤ��h_i��$g�]eؒ߰ɏ'1�\B��w�R�|2�/m��[q����\�������]1'+5m���=S������ӗ���:�� ��V�d�E $sH�p��U?kn������S�r��RQE�<}7�?����Z�#���c�u��F��Nv���L�j��K'�����cVE�6+2 ��(��t}�~�@}3���t������{��7�� �{�[��8k!l�!P�K�c���+�C�����7s^+��)��}�f��<=4���3���h~ӡS�N��r����1��d��?�E(���"=��=���a2��S�'JB��A�,1}>�V�#^&��v˯Q5;��P9E��N�ns��-̐gO�E�����N�,5��`���1ϫi��ٹ�Sٹ�_�haV��������W�7n��Ej�WU�	iM�2�]����\F�i�Ѕ�r-Qp/gdb4߶��������=6���~��NLGꉚK�}�|��ʥ H�p~�.|���)��+
Q)�!�4?5k���1���K���&2g,���f�t��}@�TR�!" �5BD�R�A����-L�;%���1J�ƀ/�����׎c����{��{��K\�H�eTţư�׾��I���RiDkp��u�ו�D��u�탧���B��F��0���_�5�Q(:.H�iu�5}L�Y���[k"�r�&}}u@M�G���O�Z���F�<�B&h�0��!��R�u�CS��ɽdz^���<�\ 
p$U�j���ڽ�K3�z��K�z[6D�h=ɪ��������o�MU�|+�Pf/���6l��9�+3�t?{;�n�suK��C�N�Ktkv;_<J��״���΀��|�@�fm1a�]/��)OC֊��7��������dq�u�@F ��~�u���4�:�@��!�\Ji�7����U=�W�����S����̝��� ƛ����ԦI�泒G}R'��KI�VmD�N/ӾVy���^X��#/w�q�n�S-�?a{No�F4*/1׿�\��QA��b�[����YC��=]��L�+���'l��*eT���m��a�~�۱[~���,Y���!m 9|����Rw35���(+�/^]�`4@6�����9��#:�R�A�kL��cg��[���d��Q��LuSn]pWy3_��SH�{:U� ��$'�~Ȇ/�@(^yQ���w����'ź6s��<L9����(qcB�(���A�&��-��,���N�bnU���j���岟�x��0�d�z�ر��r�������Bc��g�2�=0�)~Y /]X&��(��G=Է��:�L��J�=H	��13�Uk�oA~BP,�r��"%P�8�_H����*�� �Nߒ՘�t�}@�A"������(*�9EМk@�g]|�>+��U΢r�Q�� [H"'x�О��>����&��Q!a��4�AwN��G�_��ծ�c$�R1��,@��`�+d�~c��\��+?C/5}.7�t�,�6��-�u��h@���x��'Aϫז~�����3�:t1G[k�_�3J���K"D~����ܝ)YZq�Փv�&�T��v�/��y��ڜ�tD�lϡ���Wq�����C���W=/i�Ǌ��*8�i��cBfέ9)�k$���ɱ�0^w���I�peV���eG?�뎖3G��#�V�/;}�V��n�,G��.'g�X�.cX�ʦ��d���>[�BUG$����r_zN��]����[�_�˭8�^���є(� �X��R�)�rtzQ�}V5���?��Z�3|p9J���1������ys5W�,��{�%,��J�oE�FK�A�V�C�.�2���/�$x(���@��������L~ɵ�R5��"���M	B� Q�~<L�f������39��|���_�@kd�Y��$�q�EESƢs}3(�s鿗�˹�f�&�%�XYZKLF7�a��J��{��*�?+Ŧ���rܙ[��ٟ�q��y$�_�</K�W�V�xv��aP��W�����'���ü~�~��/_��������BT���w��4�i�9T6m�8�Ĺ-%��s0�6��Z{l޻�~��3&i�p��Rޠ���x���L �\^^�H�t��y�
⇜�`����Hb�b����A��r]3��c��;3���t�����?;��]G?V��?a1G�@+�gqT	r�����*Ri�^(c�L�8��Z�HK�vx�amzoX�^޻t)\�R_F�R<(Oϐ�F���2�{Z�HRh�ϪE��ޅ�r~���ET��4<�3��f������>d4�xO(H��o����ӭ>^�lV�k� :����jW�/����+��Qi�[b����l'LQ�KEp�n���L���,��{~"'T=�J�w��\��	��`���K��T�'!_0)���l���� f5�� �$��x%�b�:�Sy���G���sy^,VH��NRms�lY��+Y����{uk��k[CGN���cX���`��?�-ߙ���G,����V�2d������,�%�m|��f�Z�>��tR2�-/�(-��r&>���A>�>p�X?����8���R_��w��1L?��7 �$`Y	�5���!�+�Z�[�x��N^]?��q�/����VUM+���3������U��8�=�[�;u駟�����.)�51�}���`�@&�
]Lc�h+���)����bu��"h�2f�-�{k�"KzǷ���݂J��.k�`nB��~��K�1�z������Sb����T�_��^CO�gc�4������[�(�C�^�/׊8��(D�=�Q̈́M�Q%�;�Mlܪ��yH��x���u��xmii�k�w�c��I��A�n(�]-�)_Ⱦ�Y�<EAn��Q���1�r�Τi��o�!�7��W�l|@�On�CH�W�(]�<�}�����>�wm�߷K�tUb������ ����5K��31�4�xd�/�G�w�|��&R@�>XU��T��⦸�������9����׫���Q��uo'V{�R&Xu��_�������j�OOkŲ��kZL�2|$а�l#X|J�nf����R�@�C��?Z�d�!�Ӄ�V��P7�lo�I��E�/���g�(���g��kݳ?G�\\=d�=�������?:�����#����H治��ߩl�&����j6�Բ߷z<��wd(c�$�_�"�����8 �WK��\�}�ׂ�䱱 �D�����;�ep����^/W�����jc{r-[%��"͐l^��������r�Z�u��-��Z�!�ݲ�h���,����^�H��3װr�c�K �ᡶz�>@�/ӛ�9�}#�z1��Q��G���^Ä�J"��)��/f��*��� z",<��u2��@���z�,��IӶV�Y�������ΥHU,ʾ��J�ǃSq�j�E�j.��/Ɇ���D2��U�~xn�g�pꮮdT89��y��E��`S�:?��Y{[����#l�����������u����D��m�0w��#�ߗ3a�e���p�Kq6�(06/�x�,Ş;��Xs\66%x�QEl�fȲK�X�=����c6
��+�w~�hu����+��[+���*�MnW�0+YHL��5 O�s��tx��B��A60��HQ*�I)�%�&�EI�]_�>A�_��>-��ѝҪ����/ۢS� ��pi��&��|�&{|B����v�Z�����0'��_�{�|)��h/�B��}/�1(�@׹��$�U�7諛Ľ��R�^��z�J�%���nTr����h�]�'�;�sW��o7��@��ko����7d�� �۔�/>df����� ������8�
QF�5������ϋ5!=Q2�g~H���y��f1�q�c��d���FU�5�-MiD��h!�4T�+j���[�Pu>Q���{λ����k�De��8KI=#}hA��Z�ʎ���S��:���1
߬�8��N�y�]3�'��$I�(,�����N�O�k�I#�g�LfvF�kY�IE�Uï�E��K�2��JK7��Z"�oU�n�m(�R��",��s�jm�cl�|GY*�x~_���S9 4� K��V�"�b�Mw��C��KuN�Lj)~ ��]˿�Z<擬��&��_1��z�RQhvl�n��V���UG�)RX�y��/*�Y����4#gR�����hT�|I��F��v���k�Q!�)6�[��~h~Q�Cւ�
�ߝ48�yT�ꐀ��������2D��U��':J�YX�.�y���*bF�����k�9(�����t����k�o���tf��Լe�)��`�LR&):v� �L��d��b~h���d;���ak��9���*�P��ㆾ?G(Dq�ZQ��ʎy�*��t���Z_j�fx�������}��"!+��Gc�Wķ je��,�ݚ�����Y_�ݧu8M��9�Vڦ k@�_��� ��UCb���y^�e�ǀ]��`�7�pD��*���8;��t:�qb�$�A��~F�P�u�W��}��]`u���|��ː�_�*`M�9��i��=[���m���L>VpS��f�u"�f���k��R����:�������G��t��޷Ϟ={g�i�\
D�w���c���w���<�%�^�]g@c���;o�����4�h��$�"��ޔ�^!a7���=L�b��2��D�"���~��9#��k�&���"�-=
��@u���2��!#fW��q����u\_|g�Q���I1�j|�e�a��[^U/�ee���F�ga�����Y*��/�$��0UO����x_��0����l�i^Y�/�khj���W�G�L�`�qG\>���kE{�Rl&�r"�;�\�U�RCVb�{	�s�L�M��%���u����"���.B�w��"�������y�Q'ü�A���GE�����h��:h7�ǫ�јȋM,*�
�ĊM�.R׋��M�L�b���q�M��k��o����}V��$��WU�6ѯ���(������-��c��t��M8{��g�����r8�G4� ���kb{�<��$b��X��K��^���:���7������M�|Oe.l�D��]��g>Ј���ט�W���0ב#���J Dx�O�������T����kk���pl��7!�'oI��X�G ��3���}'pJ��,��GM̲�I�[��1����RD��0�v��S�%8SaS���N��A���4��/,O�n.ν�P=���7����A���G��K\���^x��ͺ8ԋo��1�;�Vq�ZEeke����B��B;���C�V����R�Y���s�*#�0'�_�n"NK4�6	^}s~����X�>��?۰�%�}]~L�V����d��:��f[��P����(�;�D<���P��Ŝzu�.��_C���_�4A��b���*�O7�˓��U�:~�n�h�n��_�4��({K�i���~�~9}��-Z� ���o$��А;�u��:L=R-Dg��RpŹ����_8O���$�gk~�=K�B=� �{W���}3���xn"i��^�r��i`60~�ґ�D��,����_�y
����tb
�x���	�H��;�4��&�}/��]�c�?��g4�nG�p���+E.H��Q���̣8��Q�B����%~���5�V��	(�捇�5�<�8�A-���`��`��s���cI� `���O�%�Gh��\R��"��~��߄�a;����2���D��� )"�ՠ $Ժw�M]��������޽�TT�!��L�G=�"�Ev�p[��K������XDS9�*<J����r����mM��!~��Ȅ\E���qt�	����<-�F��#Q7����]�%�/;�v����Jã�VߔOφ�u�Iء�Cd���5��;��t���\�m`5�j��P �_�=q_kZ�RW�V�l�(�Ny���x��:0���ܫ"���	6���w�����;�QBb��u�*g���Pp��b�[�L-ʼc,��w�̱)�g��a�d�Ą��fD���v�5i��@c�s�`�#*�������G?���m9$'NЌ����K��%�<��>5"�����h��s���AM�6��
�U�1�?x�I��T�t��@\���K��i֊��FhF����o�]�tZh�7���q��l{��~d;+�#*�z��:d��A�)\�$PP/T�=��حc�z�b�t�	q�yjs;%z�/{�_��YZ�h���H4-�)x�Z�԰��J_f�=V�����-�`�m�Q�5�h���?������˴�7X�9�G��x#C�ͷ�]?#�v�j��dsyh��1~5Y�rr�H�_�>�߻�*2^��4���C�J���?,���1����O��	�܍ܾ}�ε�u!��h��y�7�9��	s`�ښ�
|���N��NU�@nn[�U��U���F���[MfE���o:�,�R ��߿�o\63���D��mҷuo�F�?4L?{�A���W>k4Dn^�~hK��#�x���Vٹ`~d2�;�+6:�a,��o
�܂z��޽,ޟ�����N_S3��o�7������d���X�4��_�N�;��F8D��$����JI���ك�(9/;�O'�O�r�̦�k�+|۩{�ɖ} �q#�]��PG[�VZ�X\rn=9���U��c�a��`Q��6A9�~(���UE�fv�g�V�ʻ��Z�J�N	ފ�H��n�r�q���1��]��HL�-�&�p��e �K��Q��91s��Ĉy�'�XS�X����+䵞����WQ�0�s�#�ձ�����-��	E_�0��)r�������Q�MX1{�����������mJ?�] ��]��9oN�2;�e�ϯ�
�V�[Z4��S�)n���(�zة�g�ތp���qΥ����c�T�H�_��XuI������ց�r����߆�O�q�Qq� y�:�f��@�a�����.�T��:�2���t��z��ϴ��,>O/���הW����zl�-2��}�v9r��z�2Ƌ��֕w���ƽF�����2i���iDZ�׶���g��gk+�7��n��g5��WQZ@��j-s�Sc�o�S���}w�o�?��N���"�<� ���7)z/�_5B�{����
Wt�W�yת�#,��������v:�U�����yo����R�D��D��b� t~On��]�p�� JԩЖ�ؙ��N�Dm;s��ү���bF,����(5�&j�$w�-���R��|������#/񮰁2����Y�PJ����^Z)̟������ez(J@n�
�njw�rDcF�R)����U?���G*�-6��M!�<9����#	�;k��}�f�lk�ytu�GF32<����/Q3��o�$J5}7����b�t�����L��΅H�xk�L]?Tu�x��JϝU�H�]s�C�駽���Z	6G]ŗv;��j�k&�!y8���~z�c�V,��GN��W�@���V\�6 t����j)�����7�d��ع'?����e"%*�d.2�4/�Z��	��пa�ڧ?�6��
�>,��c�X��x^��SDۀ�������GОK?�O-�;����G�#_\z�++ػց���螾�����B��������j���@n��u����B���3Z�Y��]z;_g�MG�X�?�
/���Ǧ�TI��'F�;��iZu��f���A~�pl���o0!��*���რ�ʹ�=���Ѝ�: ړO��r���Hzk>�+/��9c~x�
)��HN�Q����}<����$G�qƈe��r��rx_�O��MF^��-�\��Nv��z��I�Ӟ�ҩ�������6�p�֫��an�Q��=���Js���F�� 8���e�28�Qڃ2V ʔ>jk�>�0�S߰���/��R-��y�#�Yk/��������k	��Y�J��Q+c~ܥ�P��Fׅ��x@rd�j�k�5�Z(X�����]�G��b}�ū�L����S߽oݑ�����GiJ�=��[���VC�LIK欇�c����\���"�����c��@zK-�]��VƧ�\Ծ�!|��g�������}�%Uc��bR&q�@�[O��Ym��~(�eb<��:�>� 8?���rzV��7ǆ�;����j\�|����g�݄)�����I�ٸ7Q��^1���SX��Cv����<��V�_a��Wn5��]�`e)�*a�a:�7�
�Oߗ�>'�%�ٶ�Q���Q�2�� ���H�.i%X��gg�>^~he�W�e{�:_h��gk����}����OG��'�HdlO��D�M諾��_���,}��3lF`~6��|$�5�K�JHۼ�,�W���c�STI51�8AƇs���T�Zq�^�Y���#l�����L�l�8]�;���Z��?��ͱy�����s�]�����({fm����q��B�{�4c�b��!�Xgd��WJ����~E'�滚��Q
d���`�Я��c�NB,'� ��i@\76:��6Q4e�?.�L:�����h�A�h�gkj���M�˭�Ϊ����nP��yڍ@M5~R�u��"i�hV�w�Q��>I{�\z�� 2�/7뮿�w8�+I�0�R'��2�~�3�'���DC�D�s��4pVֺ��Y�zv�u�D�޽/�.s#l�q�U��A���7'B.���y�#\��Ay�
�>pEofW�}�Z�'$<#���!֤��l��:Mda� ��e%�����<b��Y��e�:&���L?�w �W|�?�Z�89ë�{`���l��[�&���2s�S�*/$H�մ��xUOtx�H�l��P����}N�;���[W�������/�˗¿��O�������>���������}�C��N�w����n����W���~]�'1wF(�Aև��x���Ϩ�Bi7���ϑXŏ�KȽ���%4`x�K��O�>���w�T���u'O��s�w�^���4
2TV"�����JH��F�n�*��8��kFJ�~<�����s��q��A��>�`z���Է��dE��ʘ�;p-5��ׁ���*�ⅶa���&f<�4�YW�Y����{z3�hF�`������l���-_0I-�S&����Z!�Y|���n�c =��f��<��ի�o|�&��\����V߱�U�e��k-R9��RxG�v�W�3T	On;k.�4��)wnJ���G:i�:$���s�G~6�p��v�>V�TAXn����*[��z���aH{��#�|Go�Wo�橅2��׽�:��	�{E�W�����S;�{&�i� �N�>��8��)^�݃O�����C��~��hs�U<�,����U'��7n���su���_��E�F{:7�i41��t�a���'�;72C��rKGU��O�4��Y�g��K�����G�ޛ��d�W1�����Bs<��|�w.o�T��e~ʈ����b!�-�f�'�7�^�'�tk��V9�RD��5�窅�|q+&x�&�:���BV�@ P���M������px�HlOAj�ٗ�U������968�/2�����T�f�+����Try-AL�"�B���y�f|�Q:GMS�m�G=����{���O�n]�! �!�D>���6�וy��r��H�鯧�s0$��*��s&�Wb��R\�IJ|�}�v4�cz��S�d=��,n}iq)�I����3�?�Z����S�K@.
��L��z���a>yeL���S���K�TaL^��$��{e�g�8��7�/�:ұ�л��vϠ�,�fҢ!�����Yݸp��cև�b��̒�]��'hyT�-��:���x�W��yzk��8g�Vw_J�i{�e'��mӊ_�w�-�m#�>\8΃^ƌFAש���u�~ �l��=ʮ� ���w����CT�ϖ��������5f���%�b���=��	S$�����}�X,��X9��+#|c2� (��>y��G*�7o�?���i>��ru���s��v�@��\×����t��Ȇ�Z�=�xq��rz��n�4����j��ro�3��S�6M�B��<��#�I��L����I9��?dyE8�lZ�Ƌ�4y������ͤ��~�i��<+��=�ݩG�����S�gs'31�mdG��Ġ%{tk�HEYϛ|{�"y+G��U��i��_����e"5TZ33�+��z��?���t08�n>�3?z+��P�m��4�d糣�j�;��[�Ҹ\������<�e�a��L�L�/C��,���`i#��ݛh�r�r4v� 'Y���Y
#B�yM������U��ܼ`�R��ׁ�ڠ�n��~z�\�^!�5�/�|`V�<[`	(.?�͌�@n��Uo�j� G%������
�g:��e�k�t����7�����Y^��Y��˛H>�o��pWT�����L���@��m�� c=�y��f����7�?ݟ��Rp���ߨM���)�빅؂�Ь
���O��� �
^���*	��zh&�o|��C�k�-�4���d�H^�i�w\���� \����-�7�S����pЅQ�e�Ќ���
@.�X���沰]�2N��~�T]y�џ���{U6����-f��)���#�^�W�ڑP
��0� vcP9H��_��5���i�2=a���)nׇ�{H�a�n?�{O��k">�O�����9H_�5�7�H~����HE�N.!�j���B.��9����ku�kaM�������4��fg��;Oh�cpu�>��w�����Ɠ=� /!���ȿUS���� ��m���{���93�w{.jaC�А����3�bf�m��9�o�|cN�׵���[�o�9�t�Vo����k=s�����"kC��
�ax�*�C����0�qs`Vs]���A�J�W���Θ�1���y�Ij}�ٔX��� �?��\��Q"�딡!���Kŧo�Z���ٓ
��F^XdGRg.�2C�}O2�����D�ۦ�8�%�n4�CB"��,.����U˱{��e�M����K�u�\Qs����(�s8�Z]7�����h��9A��IQ�^a��å�eǡ� �fҖ+��Mi��&쫠��.N�!��q��o+�j��@�KC�?T�d�*�����d(���v{Xs���"��#���N�Qo���i3�rP���ϒ�땵�\SnFx�?�D��#^�L��9+�m��=����kuMcT���ӟmi=������@F�o=_0#>c���{��֎K�砕��{�B��Bn�9�Uǋ�g�ˀ�{ˇ���Q��P�����/=���N"� �y���
m\�t�#�?�U�j˺��<���0؎���M�ՑT��ĈT8�Q8���jnN4�V�X69��D�#�-��^�!Pk��>㥏�Y���S�Ae�FkR&G��3�+��C '+o��O9E����9,����+z*��GE��p��*L}`�n�.��.;��ͯ�r��)�#w��Y�d&���Ŵ
b6����mƽ\�|]����C�{,&�E-�������Cb��RTNw������܀��.�زU�|�7o�# �S;ˀ|\d�	���I�ߜz�-4�0��y�^kO�t��-F�)(�~}��Q%������`��F�>��	�`�L��F9kSX�R<��~Mc1�M>[/�R�l��NL�1l��tD�Qa����l��h�{�E0���&�a�7U¤#���_r�}����F�Z�ǚc(�K,^�.�Ut15�rK�����u�,����.b����;{n�����V�V4�rLM�Y�E�߼v�t���w)Z{Js����r$o'�в�j�\F�4�L�ZRנ�,�<�g�s�r�"��Hъ��N[���*�T��8��m6��m��*4���5=�C[$C�����
��`���)ju���x^�f�w~�����#���[�
�[�[늜�Ó�gj�ꦹtM�(Ukl���2�5%���"���`H�c��� ��Lt���B#'�ۼ����Ć޻C�FnC�63��Y��,�|Y-͝A��ڲ�.���sW����&%~�,�.���=n���t���3��g�},O`u��)=�u �����h��鮁���\����t3�&���$���eq��NLs��>|)�*�/@�LT��z�+����zO�:�*ɸ�� ��-�c��q�����3���)x��}3��zΰmM�)sL��@��:�$��s�k>�]WoŔ+c�?�ֹ��#��l�_�mc�cF�$r�v$�������K��Ň�����3�cf���_�B7�*F��Oz�T�aUO�l\:%�"{[��*�<�͂@���t(�W.`��C���"�n�=�����V��UC;c������Õ8�i*vb2�@�C7sZ��\�wt����\Y���8AI�n�����e9jQ�u���ǯ��gh�v�q֎����0�׎��8���JƆ�V&�	�:���]�������hׂ��v�;�ΫSA?�O?� ��Kj4�UA�_�(\?�ko���G���֏�SA_�a�n��U�&Q!��"�������A
���;�P�LfvǊ.�j5�^�29�����"'�0�^	��3�ۦ�"͌��
����z��'7�cnP�\�*��-M|e6wvn�['���o6�}��64��wgk�d�L��m��r/�.�� �d����t#D.�s�@�w�n.��M*^��I�^Z�%���E,�pz��Yv�*������88K��B��k�����x���=�o���C(�"���=	R��ܯ ߛ�A�G�_0p;�9�xNz�t����l<���׉t������B�ـ�w��9�Eξ��^?��ön��A篱����YZ�Z}�ZW|B?>aԥ���Y�er_$�n(��Gu�<c���;�=�q��\8��l8��?6*蛕�x�d�;m.t{(���淡R'�#���Rc�����-��}��+K�t&�E���=�9�@�Z��N�h��f�M�̪ޮJ���{���sˀ!F�Muu7]�8�!���C,�+�m-j(E~����+��9�	8{a �?�߈5�����Mo=>B=��^�&9&o-㍐o�h��v��mTW�[!�Y��J��Z�S�И�-S�z�zM}"�mGA�"��S�|�U0��`�'�V`*R�&Y�ZTZ�ʶ�Ki����,G$ZG�ϔk���1������X`�;���	<g�<�u�U������.��Ž�>��Zt.Í~���v���^�����fg=9
nwe�ʖy<�wo}Ѿ���uW�W��l*�S�*0�����z��@���L�tH�p�}�V%��䩍z���0�z�D��]�W�86 N� ,�T��(�?�� ��Dz*II��c����`�#Y���
(�de���(��8�U#+]�L���K��)���B]��BTZ����l�E������L�]9��^�r�wޙ����'j��c��v?��$Uf��N�#)u˟rBt��XX	�j�0����c!���&�R�\��F�9�sb����b�P�W>�Cf��tF�� ��A~�tL� �
�lS[�Y%��3�bN?Wvߢ���1O��#�����+�S��Ϯ�E?��N�^����5�Cy���i����H�Q���\�M�(ejϸ��X.-�qЃ�L5��~����a����n(�[��]��H�;�7���+�0��_�����Ë�����b���$ yIN�0]v����_��R����RC�z���	�U�l��G8eF#I��g��_%ꋮYD�Lʽ�]�Τ�|O�	5֯5ddf����Ȁ�G�-��l��Vl�BM���]}�r<<��)�<�Ϻ��Z�\�_�H9Ʒ�~��=_ëk��P����oBd�[+R=�@	��_)��#,�҃������c�\7�;͇Z�%�<ZRa>D���\�(�)KI�8�8S���>��U�h�(�s�ޛ�?a�5���W	�cD�U-<}c��Fm䤑�jv~8��L/�%?T|���tQ�s��E-�S�`8��\g�s5<8��;��O�-�1����ޥ;F�Y�dȠ,s�p.+>B�]}�f�S�nY�=�ߡ���3���=�n�������W��������v���+��?Gl%�_K�fy������nZzRW[qW󮪕�����O�;7^ap�Ɔ�Ez+�9ܱ�̋Pm���b5�:5�h�lV�Mj���� ��~��7]�DE����_Ҭx�Fm��3��6���8f��z�`����.2+c��n�_e�h����X:=q<K|��f���B^��y�	'G�	��e2k"�j�~�7��ȉ�&��}ސ	!�2��|fw}u#:��K�^b��`t��2~��X��0�m��5�$��f�#׍wF�6X2_)�)��5��ݒnBx�ԅ���"���rZ&g> ן\���[�]���@\�xZ!iˬ�4կԨY2_��,7�e��tn�N�_&;+�T?�l-��g��Lu�Gމ¨���r9���{���#1K�g� �W���U?�Ẋ�x���N�Ɨ��2Y��'�����̇�����e����r��
�l�aX�����"�@�N(9o�
徇��Q�$�^�V�Y7��j���9���6�녏65 r'҉@�lqő�l�i���=���zM�r�)���u�Hި�޿q��&LS�'��%�t�c�b�H6��U��%!b6c���$�A���������#�n"4o���h
�s�����C�ǣ
�A�V�-}��)ꚰ;3r����T�p�t�oO���!{����b�{MH4�g��}�iE:<��n��Bz��f�G��[���<�c�<"���L�Ƀ��._1ug�%|h� �7���,���V��
sGc�5���D�W�MW3�KY4��ϊ�ω�/��5DU���i�	�x�R�~�El�A���X�K v�ݡ��\c64�J��#BϪɻ�͑�[�a�9gS�Y�j�5'�_i��%T�j_0����;���]�|	\�F��1m`<<Q��>#lA��/s��M��w��D�U��'܂�݌{ɳ������3�ue���?B�`r�=��(�,��M�N}���m��E�vr�39�[`�鋿��iX�(xb&�۴9t��ʃ�dZY9HT)7�Fd�D�	^~h��^�2O�Y�W"7�P�=�x���CP�h30U�1���D! A��x��&���D�VPsmAq�!\��9YG�: ���J3M2���]�γ<ZwZ����Q�a6LG]�����j�^F��{��W��g11T)i�B�Zu&x�������k+��B�$��✧v%n�q�+�Ag���}�}kh�J�޹l���eMb�<ڀ�gp���{0�7�p�!Xۏ��u��y��@�az?�/&t�	�R�zS3G���@�`��8f\��BAVs��=w�lDk)��=���b��!�[�	�.���:����B�!���g7BM�keLK��ʟ�.�Q
r����g�|.]�?����kJ�G4EX�J-�u�x;>����V�=�����ş�/�m�n��⧭_���jF�s����I��- �%��Z�a$}x"�$>DB+c%��
5�b�<����9<����Pɤ�.��{S�m<Y���OP��8Q�}�g�"?Ν���8�鰤�"�W�.B���R>��A��2uo��q�aU�:�~�=�O�_c�F.�;?R����(�e*�l��cmַ6'��aA���]s�5��ܴc�&���[��r�����9����]N�`���|�ʍ>v�BM{CE���Hu_�D��q+Vw���(��^e��l`'^�&�Ά�/�E�s�F�]Ѽ�ӽe;�b�9$��x�m�>�8�D�`�U�ɩ%�Π����\��|��\���{_�ap�,����W�p�������jf���U�{@�_�R�S��2��$��Ֆ��L�Ƣ�)R)(iDDh.�hN��(%�ru�Uͣ�<�/N����\���8o|��gHjv�:�.���� F�$��k�L�
�g!]���h��Gp}��li�f���B�{@�ً{�%7|K�Wn��q�=�\�k����w��Pc]��j? ���q4�V��r��CGZe�f]l��۾�[/��a��|O��k1?Iނ//�9�%��#��wF"��Y���ތ�\��d6#2~
�}������E��������ɑ��9���緹H�W^!�Q�#F��Y�ȧ���>Sy��×hW��c�s��&�8�iG���B���K�����a���$���e�֬zA	7�%q<E��-��������e��e��5�yg�F���gp���ƽo���:�l�d�������ׂ�+�1�z��2&�#^edMU��98<$!X������k
��%�@����!���*��ʎ��5� �M ��[�m�e?^���w=R�c���u�R�gt��
c�b{K9;Xy�%�[�:����33Ӥ�S���]]D��Ybj��Ůl눨gm,��~��:ɟ?�q洟��<h��|��W��|��lb�6 �Y�������=����F�D�� �DV��K�ؘ�
�F��/֒$�" -v��L;ԡ0f�L>8����72v�]�~+N��"L;���T�&YF�O?z�;��$s{ׂ�1c�9?\��|��e������fi)�������������������da?(���m<��ss֤ab��5;�X�׉�MBj�MoTj����q�w	�ZJ�V"�sS	ѧq�9L�E8����;@�U�A�k.���Ry�֚�A�6��
��w����.���Ը��\�k�.a�E>��?��c�-EBi׻�����ݳ�g8��'*��&�=�cv]�<T�h�E���:Ts�ϗt����U�ܷɶΚ��Lrʎ8�Km���S���G�[�E�F4R�t#�R"�t�t7��-%�C���PCJ�0H� g�����ι�����yb�{��^���tY�?�[7�'-W�lK��d;߾U�od����N8�����5#�������0k�߾k�D2�=:�-��@�\�ݧ%������z2����4X����{}��x���=�O���
�^��ē�����T���OL:tk������_��ȋb�?��Jz��� �v�� ֐���xݙkC�(!v��0�;8qu��7���ۍf_C�s=6s]����6�۵��%�@OFe����m��A|2Y��\�`�����k�����q�?�j��/0�:�y �������d5F�1^�*��%���r>��>�ڴ m�i[]�~'P���}1����o�8t��ʘXݖ�}�
���w�.�̌�y��X��>�nB�>y�k����
���il4Q�ܮc��]�@)�b�Ob.UOr�~}#-�Zn��9����LFd1�G|����� �X�L0�	�<d���5{���V���0��,���,�]+D-�\u4>墢�;�^}Z��`�K����~,�SA��f2{K_���$��X��J:���l�֓�o�N�(F8��8^�_P6W�C`�ZeF��9o�&򮁤mз[���jKX߉R �)����FJu�M�6<{E���N�<G'����Jͤ|r��X�KI�����ĺ�����bd\���GOǔ`9�f!8�^���2�S�-�n�0��(4�:���v%3A�ͯ��XL9x��N���f@|��T6B�?�����a7ɐ�}{�� �������|ƺYz�K�W�ND�;�c�s��eQ�k�g*��o:��44V**[��^a?^�`�W��f����F�l����d���,��θ�o�y5un^�Rw�f�k�1����5��ix�������q�E�\�G���
����@��s�0G���*�H�4!!�,i��i-�1P�R{t�����Qv�M�6Z�s�@�%���,봲�W�#x�g���Wt��J�'�A�`(es��M��<��>��\?��[�ݢW8z���Z�����xc�%�7*���ʨ^�Yz��KGa��5L�G��T������O�,
�'2X�'J�|~�a��k�p���^��"E��R��Lz�d.� ����c�䢸q1ԊA���h]�?~���-�5w�̩��N�v.@��2_݃� Z_��`K�������@Q��I�}�:t�/f}�f�,�h"�.�c`��k�n����V�LF}{���MȱJPUE'�Yܶ�Y�QDe'��ͧu�@�8Y����5OE�ZjfyuY��`r�����}��a0p�r/y��Ɣ3L��?�T�p�XʤH�m7������o�?q�o�������cb A�Z�Z5T7	L�(auB%�2ջ�q�E	����%.�:Q�1j���K��tJ
���qh�ֈo�/���+�$�}�����W���I`��a�M�g��:G-�%�O?=�]:R��?�jE-<�r��4�����u�r��J�'�	��7��]���)����(;R�o��Q���.�w�]��c����u���*E�߉0������L�U~�j�tg�{����j''���Tœ3}��@#�Gph�e{v�[_챛�@�����N�a��~�Y�Qt�ܙ�?�N�����*���@�$,�]+��J:�������sԫ��'�R�����o~a\.�Û��� 1ɠ����C9� ��b�3f�!�~�L�?��˖rny�1<˖�N��N��@'�]v�	��bB��5�n!�̶�Ȧ/��a� ���de��vbk��Jz����x\.y������vPPr�̆W�7:�)դ�	���NJ~u�j)�HY��0B'���_l�������7|=������^�Vk������B|�x�Qmt���K�A���uf�{3>Ѥ��7<2���x��妓u�������f��>�K`�,G��x�P�\��\2��8��]s��Pב�$�I5J@s��ܲ.{�
mlN����ʐ:�EW(�&����$�A��JG/�&lxF��
ΠCZ-Er�.��H��]�0�ELӴ(Є0'7\��Պ�{;� ��$ԋ˫0���4嗝�vla�q��p��ּxw�ծ������peP핋-d�	���ב��CCV���礽9k�k�fK�{	|4�>���nς�?��0ґ5��Z�$�:A�`���?Y��Ș���6��V��G��#O�ƾ6������\�y��>�8�d4���4�"A0:�,��u�����cLm=˝�.�Hs�E����1.� �8�3��B�U�c�B��?d9fܙ��P��C	K��Vմ9�	�n��b�Q/��bu9{u�$�q�E��κM/l�%�昑���8L�q#S^�?
!$�m0K��ɿ��$a}�j3�]��	�
,�>B�J����:Y� iwUS �t�Z�u[�-���S�Y#�~�!;/�z���.�eI�4(l��G�;�>�W�����4�[}	n}�;%��O$}h�f���v=�F_�o��"��o��3��.��,�K�lW}�J����_# ��nQ�83	3�����":io;�d�,Ҍ�c?� K��	?Uޘ�)�����w����5o �dh���Ϙ�ZA/�r.M����f������a�KQaݟ���U&�V�0�����ʠ�^�t�-Q���Z�bnk��4�w��OI���$n���]s/T�l�ۦ���>^eP�K�_Dyn���rD���.�˴�G���ݭ��?�!b!馎���x�k�'G9�䚚b}k6f�r�
&;.R
�����z7�oyӗ�~k0Gs����@����B��>R���)�OJZ9�їw�"�"�m�g�s��?���p����|B�T�j�Uo��?�R&m��'o>��0\��a�R@F��t�c�==�L]>Se���f��?9<a�+&dV�ҬTE��A����'�>�iĶd-o͌=
�㫖���~��v�b��c�;ݨ��ʹ��k4S����*v�9�J�;���3g�]�f�<'s	�5�2���V��CM��S3�Yj�6��:;�S��y�B��c/��n��l�ڶ/��g���#'�}���Oz��GdG�y���^��C�pw$��!����-	�݅�,���+A�=�񲯮>`�uR����ol����0����*��� c��?nӲl���oKs?ƨ'�A�N\�y�N�楯��ڢ?K8\�/������\ν�a'���p��D���c��
�t"��������DD�CW����_f�V䊠�7�ɻ��yGu&���/࢛�v���ڐw�B��Dǡ�r\!�.�S�;�8U11�'�Qn������1�ڴ���������0��%�]���6��Y0tP����$�U1v�/�|k�t�y���l��;_�����YaA�B�B�s������46�ިT�Ԗ�Kԩ5����;"�Q��4�ގ�	�����`�S{���\�Z(H_6kа��~]Y�޵T>�~�a�~���CLZĀ���ք�,f�K(
<[���[��}R.�9$ݔ:Ag(������"�]D�-E2����+��u���Q�DE#Q�T"�xզ�E��o�D������Լk^�\���ͧ�OO(�hnWpܢMtI��py�D��#����� 2I��T�?i���T)P3">���J���k��;� "�LfW982��/㧹
*�M�^	�j�!P.p�N�2k�gQ�˛ +C�}]�E�2z����=ȉ�w�Kr��U�e�8��4��4j^�#d�1�Zc,�=[���˻�����P�`�_$�Fo��N����Q>M�"�<�����1��?]U�M/<�H�M��[b�6��4���n�
�\b���L�5�����]�29�9�Z�O!����}�q�_�D���mn��{v����Q�W�Z�%��l\{ηд�s6w��5�,ۤ˖��4渭ʳ� ډ�]�c/J+u�� �h�	m��00���쎘E�b�xF�s��� R�#<J/h��_'�GN�e x<R��%�C���je�R�3o����;�B�Spe�׮�2�<xh�$�	ʡ��
r۴G��L�����z��uJu4a]v�Êv&i�[�$�wL�2'%'ۮr$e\����ٱ�0$百�V��>��˼�0��tZ��3�����~w�f�s�L� R�7�%`���-�Kv�O�8��8J8�/ũ<Z������U��>�;*������U�����<�ϱ�������{ٿC\�Ez;�}�t�J�M��<�$�²��< ft�����Q�F�o$�W��BF��Ve�ҝᬡA�y^�^S�y3Q�rc�Y��g���$2+�������:��5��@�NL�[�Cg��<�[��ˌ��(=�r���E��iM��{^��A���aw9�^���㩇C�����?l�"��I�,�p_yP�k�λ2V�{�m,��G���G�Y��Ῑ���w��X��ʄn��*m���\�����G��\��7zխ�5���f�����vӫ���b���m�
����Hx��}W$w�:0�=��q�'��/P�n�F}����57�Tn����c������^M��>]^��l�c��9j��e�/@%Jhr�$�Qm�=�8�ۙ�}w� 29m$ rKE��a~�W��8��Y'㵜��h�����_6�T�K�!^rr�(sQ��|o'm�[y�o�۾3�䒗�&>oG9M(*҂����9;��v\:��E��p�߇uOo��,�i��X!&}m�~W��y"��+�����@�9G֥۝����8`D�_���h���5�+*bp����䒕��܁⺘μ�hUt|q�r5PV�'19X�7b�FA����:|3נ�l�l{�D�&
�JD�Zw2QW�:ѫ�����L��̿�a�8|k��g��������H_����oQ��W�Wm\�r��UP��hCC�/�T 'P�y�7�}�ϲ�CN�-	U�Z�`�V����l���t���M���L-k~�v�5b��B�(���=+�z`��|+I��[��rB�r��.y�_�#u�֒a\��r����ǠJ��c|�z��X2����r�^�nsړ\����Z��/��fɵ{�{Q6300�B�:�z�y4_�=vZ�����ߧ�꺃�_���,��ʹ	��.�JJI��� ����4I������u�r:JY��{;�
/�=����x����A�����"��؟y��s�u?F��u�ݘP�������a����aׅ�����d�`U�?~�SDh`pW\��z�D��_���S']������s�J�5���Fw⺸�����&,�]d�W�E����=��	�㤖����hs����vlҸB�o�Y�V��޳���C�!�H�������=��� ���6��f+�z�K��ӄ�L��}>p��d�sU��+�0h�����gڳ�`��@�_��X����"~������eVx8�(���v�ɏP�|?m&��7�pB�ɬD���q ��T�hXN|�MZ��oo�{S�I-0�uf��YhtNt�
�5͂f�|�������輟
�=���v��[�:�)�j��ï_"e~wX� ��q�S�z������2��i�)�8�R-K@�㰔�3�����@h�ڸ���{Rb�w~/�.m��J���b�t���8&֔��e�T$S��X��a,������1������ِ��b#UZ�	�o������PW��!mkxM���(�i#�9�V6�T�+B����o�ւ:)d
 ��q2�CFʾR��u����.��zy�?�`�{ĴN�<��p�3?6	zȎ�d���0U��,"�wzF�����fL�e4L��	������0��hz���k�'�pL�䒍,�M_!�Pb�)� �i��y�J��5�%�ȐJ�p��=_��f�)�s�ƹ�^r�顷R�A������6�`���',�>���
�ol�������Uh_���Ю��G��>��-��I�����u�zS���Y����l�r�U�*Iq�ݲML%<��b|:O^f���0��	�O
�W�?����]G}�5���|ׇg�%�9�^_�z�+�(�a�8_��t�����捐�u�R�Ǩ�_�dha�=CDK�I�zƣֹ������ƻ��x����{�Gc!���i��]L��B��<���d��2q����ɰ*3��ܛ��7��{Z̈t��pp�@Mhe��z�6p,b>��tb
������H¶�K��L��qo�;M?�l�QP���!�뛣g�x�d����S\�q���t��K����V��'��q�ƫ��ٴ�SS��VM�`d@�UY?\P��K4���llHo�Ã/'�	z5����SyZY�'Rƿ�n��X�:�m�_o��M���
���'�21����۲̧q}�P��g`,�Ź�&���ȚT��Π�|��Pz��"}�~"S�.a���<z8�2,��z���y�D�7�|�������W��<佰s�g� ڧghJH>-�����7D���G�{����*Mzߌ��Rj߀3x�)bbT�Ҥ�?<Vpc���bn	�o}s�S�~�By����5�>w���N�� ��V'u�y3]_w"��S�{v\m��}���W��|�8���v��V0���$��V诂�6��nӧu�|�TzR���+���þ��3`��X�\�][Suw�°�u�*b��$� ��j���&4[e&!)1�iw�FAK��2�@ݟ������WY�
����Q#��`��
���o�ȑ���"V�֬b��f�h��3���jp�oNbl2���P��f�Hd}���9,���X~�VH�vQ�*�p��dI�[�14�E�
\|���̀A^�~$b
]F��9�ӄ��;:�z�{$�Z������/�>�%��f�~T�v�.pk�s����������;Ru�t��� �H�D
r��bM�'`�X���j�a�b3�H�������H`�Ԁ�f֛�]�m�'AG�	�ܪƎ;R\��&8��	mK�"dR�}�Fi�9��l��9hhY����x��$����eصgȸ���ֲH7z�Y %)���/���2��MV_��4.�1IR�n��݇��c���r�1a��T|z�b���?����e�p�b��8p��dƙ��~%u�J�d{�^~M�\��i�[�O�X����&Mc��݆���s��6�̀��Z��;��[�	_|�����k-W��J{7�ـ=z�v/F�c
xb6��÷՝9,?��螞�i���,ͅ��f@>HI�{��QA�����#8�q�˾�A�v^�����X"����V�^�;|��J��Y���������R%ܕ_����]�m�I[���X��{t��W3���4�����;:�k�}�m��޵W^~��~B�6��CT�^�݄A
p��`ߵ�;m�(�Ҿ� �|�����.� ��Tll�k��w����0I�!d�;!raY�`/ }��  +p �qv/Q�U����������a;�4�J?Z�P|��w��Z��h��7wZ�D�EVj�^���7�XW��PE2��	�.�+��5��E��n�s�l���z�f��w���gX��X._،��*�gy��������x��i�
�N�q�}4V>�L��àlM�T^�ӓ,=S���&a7i�U4k�O}�sF�qi:Ŗ>w@G4��`ߧ����&s�g�����
@����
�G�v�4o�dᇮ�$� )H��5-t�>�{@_`��ECG\�w��z|�.kR�2���!B2�}�S��c��T�V͈@G���ܹ�3P���"�^�E)^r��h�5�h�^���`�n*kq���D�)�x�^���rS��i���^DH�DLN>��՛Q{�6،������'Å��w߁��~�/���=��pP*K`\��Ԏ��G�=h���Sy���s}�ۆX���߂Ƚ"J�#�ڗ(�P�_u��c�@ᵼWW�G	�_�z������%����;B�%8��q	�&�Q���E�`i;=妣ثgA7�����yW%��!Y��ll��Yog�5�Z��.�A�]��u���8<��Dt����;����/��O(�;~�ߦ�&H9>��q�2h�>S�vw�{����j`�Ɉ2�e��h�8.un=
/��b�dG7��I�74E#E��o�5�GTh��h��w�g��'mxZ)�:�o-�V�d���_����ktV}��e{Q�U�Ȓ�mcB��[�AS�q'M�}���43,Q���"S@C/��C��C1	�ɴ��E�KZU��h�["ģ�����ؙ��h���G=Qb�l�VkWD�/C��S�Zj����DN��:�.^'rB�dGr�PVEq"審c�fج�(a9[_����4U ����I�L�`�ک�`�'_B���oEr���V4@��[�Bl�E�����k�x
�g՘njq��U5�lA�s1��J>������I��˶f���f��`i��p�=��os��r����ٚ�B��שY���Kݏ�J/n��%��O�cn����*�VG�̍o������q&~�N^��k���L����љ�=�4bђ�~q^l���1~цu�1w,!�c H�R	A��)X�AYƽf_��ċU�(ϼ����^A�{JH�.k��m��N�:��ʀ�q�{����s�G�~�ڻ@�lĮB+0��l����ez��K�����B�&�Gq���Uf��"���e��'��q��d����.TQ�\Dg�a�b澎�n�2�����e����ww��e%��f۵+-^a����c{z��ʷ��+�M�9Fbjw�[pNkp����
�z"�K2��W�1׻����������j��L[o����.?�}D��flBi����F(P����oh-,�,�� ���\l6eY �'��$�3"�����E]h�bt��ʊu���O�l�Q��H��u�_{����gR���mc�:lH�7�RQ}�5{�^Ɵ�
z��o'�|��T��9Z�L��V5D��6�����U1��J���mp�Ủ�v��Qi��ŧ�� 7�ҷ5�z�����M�����MN���"�/��A�)?g9Or�v7U_z~��ށ�L~ɼE��A M1v:ϑ-��T	k�����T��r���+�,5;��@�"���:�>ͺeޘi�\�����ǵ�$k��a0�;�	]y_�Ch�/󸧵�>������������0��k]�O�l�Q
�i^H��;�ߒN�
5U��V*�kt+y�	�����Ч�쐍<ӗ�|ԁ,ݖ7�0�j��e:�hy�
G�޲w�VUݕ�Pq����h���2.A��Q�d\-�H	�%�s5.��� �~� �<n�˾Z&�> >7�<#JU��+�3��R�!BЮ�$8V1����<+���;����fx][����d�[�|q�YK+�	�c� 2�wNu��il��E��N[k����8��v�7��L1���tc���2*h:��UR�W�O�lg��h"2h�D�G�3WT!�w&����M��iV�2Y��'�g<��dNa�T��˦��-6������b���]X�<�s��o����HT?t�k�\�S\�x6Et�;N�����W���록ڪ�^c$޻.��BvG�W�Sk���r��ݔ��Enx<^W.��y�3o�H3�<SL������ -�h�0�ΐz�/�GU���?��lx��1�Vf.ϥЙD]E�O�J��ܵۓ̞��˄�f�������%����o���Z{�W�;�h!���d�[�����z�Z;�#	l7T���D�	���y�H .�:�L��}V804aܡ�Νe��x�mI��ӼꉙI��,����s�O�s/�FS�q��T �G�&(���Zs?��l��Vv�g=M��|(��b+.@r�S��ۣ�����`B0_.n#4��{;��޻�tB�����&�nwg�t�X3YZ!��=m4Ua m�ҁ,��ơ�)sQ	�5;IG�	8��1:�������m��޾��HcȬ'0�[Y\ޏ�����˗�T�q�����Q3��=f�5n��� O���ӟ~������A1<���+B/騒�빉�2b*z� �YQյK�@_��$���K)��`�p�_���;�>~����(\'���ZF��;Cq���|w��)ۗV�l���e��s]���M�o�,h�� 1�$�v��2`[Y�s�l���JMx�"�?��f�s��D��b"gsN%�=N���{pۻ_�-Ww��N��"�kH�Lcd�T�-�W�Æy��O�Z�P�."�9��1��,6~��߽`�h h%t�WWk	Ri�t������0K��4�
�caҒ[#\��s?������nς<0���@�ѲBKX�҂)
���Ѩ�bPM����U�b�3�������x�I�:g�g1��c38H�> �o����]O�����tzY��FˊT����?rM�)���ڭ�4��:r�u������!ͮ����g�~NB��c�wrE���^?y�,Ӄ��.o����#���y�Q��� m��hG?�Y�7�� H��ddy�x@���DX_kB�+�i��Ջ���&�*���C�sD���ז��o<��Z*�ڳ�O>D��[�%�)� %��'��?$W�CFK���n�_�]$���8����G�R�1϶{-�lxkm  y�}6�8e��Utc2"��ٗYC�da�yGs���@�ɋ������t�m����s`��ho����6�k�^u�r%�յ~G�@���vIO�ygo���9�IA?��)+T�{�l�mt��b�B�B߹ +"�t�:�[�Lm7��07��[�f���i��揭�Y��"z(B�O'�~�
�#H:�G;��n��ȸ:�@팡�m���K�;6�+�nS��w���6�!�6���n��q'���/Տ���lS1)��jߧ��qC�Y�mGd�O7ҥe�� E��T۾}/�tm,�W�I���x�.7L���
��<��v�B����^�~�ׯ�ᨚԌeh����W����x�ygՏ�'���!�5;sf���|x���N�~�wy>T�(Ty���v��{6��c�'�����P��jJ�T�������_�n��x+5苑GL���$W�I�����Q�ˇ�KG��D����l��LtO�<t�Qgw{�1�}���<���*�_��8�+G���%yL[����B������_�Ť�9Q������,�1Ş�b�
(F�J���e����l�<m�ņ!&Я���.v���no���qɆ�"ZQU$�t�D}#�Q��bk%p��n<�}���z۝@=�&�<��&Vc�_#�N�"G�^a8O����,[|g.�ӧ;M�JsZ����RpE���4�}��A ��$��(�%�or=�'�bA�v�/�'fӼÖ%6�m����.�yE�}U`�zT�����nPL(�s�Vf;<k�!�V�}Q�P<p��1�U��5V$�D�	?@��'l��|g��;MR �v�C���������^��smb�\�9��ؘ�������R�z΍��dC�c�c�E:)�h_���.iE��7R'-Wx6�c"	?p��A����#$* ��9��+�zLhKu��%���=C��Lj�)6�o0�ElnDgeS+��p��ZS���]�u���4����Q�Yb�������D=�)����HD��Y4�F�]�Kv4L�Es5�!����5���W�^	償��/l7�U7]�O]�u݄�b����P��3�4OK8�z`N
B�9���\�}&��	���&=�GX�T��%�͒&�J�A�A�N�:�В ��p��K��!��H=,�BmVʇ���Ӛ�ɚo�+
'\<�͆���r��͠�k�>�ם՛'$c}î���[kю6h��Y덄U�.�{�Ba&ӝ���C��@�q�����]�K�4�}��|C�@����<*��F`Op�;���ʕ� ˍK�nc;s�I̒d���*L��?�l���?Jw~�KF�h�ux�ұ�F�k�WFӀa|*=���YU�?�u�4b��ec�J���q���V����j�E\�r�i�|��3�ފ�j�i 0�Es��[�~z��r������P6��Y�,"�m���Ǫ�'�O���`V6#��6�t��O��4��{�s�*"�YCH�m/|�����U��o��'�s��ۚ�K(�F+]\3�}�.���q�Z�����0l_iӜ����Ϳ��;\_�R�?^Dj�C7�Xͣ����nΒ��D��� DS�l\p���h���r�W"�}���+�I#SGj�b��lP�A�7�1$H�] -ߺ8�:�Zŭ�� t�H��P:?Y`��_�����HJb�=�1���D�W��A9��RP9�&��-u#g2�Mι��U��mM�~ߑ;
�}�X5���{Qe:��}4f����d���Ǝ5�M�e6������OQvDn'�
�${�<�#�&m�ݘ��c��Û�q/{��v�$�}1�=΍>j[�IB6�p�#ls׊����/SJ<�ڨ��W�|r\iL���;��yN�`2qq�f�>+���ei\=�����~���ټ6iD#Z�D-]a9�I������^GsD;R.F�Yʼv���?7
��:i��c];9�#G�9[���%z3�v��	��^2�B����b�����@=�z-��X�>����*�7B�<���֩]������J�?mw���3�h�D�y���b�=���v������^ !j��C�LX����L�3h���e�
� �KD��C��EO�G��P��4؅�
�K��b�jr�V���mP��r�k����rG����U�+����ާF���Y����e3��LH߰�b��p׻*U��f��}�W�E�b�OI�!�vɴ�.�H��*��n	�
�[��DM�lv��ʾE��T�����3��.�j���	b��/G�Ѵ�U�����h��Fg�ſ���/V��p�@�7B���G��3�57�"C�ϜG���o
����>��k�Z(j�iw�ޯ� ��=$%�eXY����]���,�����O�}��_��B[��g��5xˋ��g<�/a?ٮ�����2B��6��L+����ԉ9���$�'���jzd���2�^�o��7�Hv�������PN8�2����O;�<_4�s���ˣ�^Y��fZh�oVO�>��~�}�Y؋3��m�r�c#�߾�g����C�G��5�nI0G�i!���<�[�>��O�e��~z��!��wŊ�Fzp�=|�.��#��@@&���:a�̦��/%��gg���R܇� ��2 ߧ:�����Y��>��[N��q�Q��xU���g��t� �-Gow���L(��j:@��r��ͺ��@X�#��%p�/ 'Wn%ߞ%�9�ڜH��:���$t��bZ/�Y"�~�Tsoi� N�Gzk�	�Sz��x۹,*n`N�R����9�����?7��<�"��dZ��W�ur���uj?���Ozu���Pgu�67�����X��#{M�����]�,H�����s����-�9ּe���_<��Km+f� ���\B���蘏Jy-�3�=o��m�n+<\xυț���x�L*ws�C&�E9����	�y6}�X����%��4޽G�D��fn�p2������II��k:'�nĔ,.q�ޅ�5�>��i0�W��\�i���C�St��g}K>���X--	�Kƍ�4�F�ϭ~�i�u�H��b��Đ���p���M<�d��(w��T�*���
������'�`펍?��b��g��K�g���u�ʹ�g��px�VD��4��sw8c>��E�ȏ��i/�_<˷�-*���oLL��Pn�5��������"&tJ(~��Z�&'��Y�)�
�5i�m�[ks���3A�����f����(��ͣ��O\����9������ˌ�D5dE"UC(U��o�K�'�/�3�;E�!���G�З@I�!`6%8�˟M{�j�?�~���yݯ}v*���|�P= �^BUAᲈ�jl����i��٠�pl��67���K9v�E�z��=�_s&��o�Hn+���*��0X������I_��9�Il<k���Z�+̣��r��*;��:��[D�yU]88G$Ҝ-�̟<v���|(e�t!�����k���h(и�3^��t�A��;�������3<tW�{1��_�-���3+���3"Í�v+�Qi}1W)fq�ԕ�jH������<4W�����X �Ho�����.���Y���|Ion����+�W���[�c�ǁ���o�n�vR��:Y�-&O- 8P�/^м�G�X�d}NT���1}�l����l�,�dC��X(%�w1oEI҇�^��R;�9��;K�)�d�3�Ox��y��o�\�u/�rO�ڌiDmk���RA�G�n�t�����>�>>_���lR��:�y��Jխ��0�&������ӟ�[��g��v�7��56�e�>W�'�;T��ƶڤ���;�:9����͑Թ��8[L}�#�p�ź2F��� ����6���y��N�������:Z��L���篐�kN�i���$օ�1�t~�^>|��J��y��B���JZ~;�7)���֯n�����k5��^�sx�"!�}���l�B��XM e�b���k�cB���%4��D������2����;݂	,{�b3����,oq����?,�<k�[`�2�Z�8��^�������Ô��0j@���o���nc�q}�i1|��&Bh��$�6��?���r������[S���P#�?!���%L�^=<��?3�^:t˒@�M;>)1�.}�,x�� ��(
ڂ�&��Bڲr$v3%x\���J�z>���l�Q8k!��i�8��Ѿ#0�S�ѿ�M4N;4�,�t�p�h�E�OuNpҢS�O���N����r#�v��nܿočS��!;~��
dJ����"Z���=�4!D�ż}�#���UN��M�T�(�^:��<�e]�JN�6���^ܑ�O[�n�4�L`�1�)��c1N�����BQ[K��:�E��l7�[�C�^��B�{�*/�\8�~u-��������S���v��k���3s��x��`ށN�ىb��1��J/\��I��E	�3�����K=b�y8�Y]����
�����T��?���U�����'࡯�A����ck��u����`�ں�af��C`o�lG�%�P +��@/�#L;mUol-S;�Ĝ��i4�8�&g���@��U�V"�=���,⛠oĎ�B� ��pʦ76콈͢0R����b�E�9���6�Lk�z����A��(��~F�ӓ��Zh�.�����wtr����%r!%#����4~�G%�d5OMe\�;���R9C�W~o�?�JqI�{�O�z��e� 9�}��'����	�<�m���p9e_x6�RM7�3|�5acR�ְۢgK�Y�ybAD�r� �t��Ϗ�Qf����L��@�����<H���ߧ�PM��j�V���9��@K��D$�n��'��ô�f�M��*D1�0u򜧶z�o�.L���b�	կ}m*~�ynw3�ͦ�?�%k���7mץ��cL�_��_��w]�:NT8��v&��-�^OaSA�ܢ�z�P����C��1��U¥�֊_�J� u�����Sq]��f����S�7 �죹�~�Oz����ʚ/&��R ��q?�η=��i��ᙅ�fZ"���Ltx���)�K�`)�D�Ɨ��WT�g�ç'7������}R��r,o�����8�p����%��{��R7�w=���Z�i����Fv�F�ِ�r�i0zU7�To|F��������s'��$�yi��O�������5x��T���[��f)��_�T>mn�[��6�%���x�IPɁ��^��F8OM�'�L/�#��B�����a����2��yk��x�|0��YKR;��a��S����GC��}.�@hp��:���G��A�g�w�_�0|f6>c��	ѯK�g\�.��K�d�I8[V��}q�����^���`m��B�f.4�}�Ƞ�E�s
�2�1~W��i�?k׀L�KC��7���`CLF���t����n�ͧ�mv�K�>��o�ړ ����q�l�Q��T�'�-^�����܊�D�m-6Q'�9��U��q�:�8�g3����l/��E�9M=�n����oL7���Z絽��"�Dt?Im?��d@ܷ�$�`�7�l�T%�p�q��sz����p���VmK-~��/u�uS�|��E9�����7N�ߏ��R�(�.__I~���{��Wߘ�r��h*uK�<K�y�d]E�P�Rf�z����U�X�9����1^�[�����H*'��{@�}�u�+��5+���?���[�z6.|��z�&��xA7ҍ ))�J�(�"  0�{�H�HIH3�����0:G���{�g����}�s>q�X����L_M�yq����}r����:���M�&������[O�I�!_����K`)j�s�^�?\�O3����g[��7��ۈ6b�zA�t��83vS�%&�F���>1O¥?�b��M*�UC��A�m�9ci��g�x��!7�-0(�PJ�UD��l}����l*A2{=w=E��B�s�����NQ�)�7���v�I�9>���<I�^�`��ՒX���d��"X�<%��>����u?�N
5�Z��ϵ��s�k[�A� *���2|�i�La����ݥz������TRÓ��9�kǎEpe��N#��z�oٗ���[�lH��<�7�|_�	�k�9�����'�%\�*V��"1�'��Ac,�"�3�Z,&�e�'3�K·ؐM3	�ɹ@ܕ��:����UU��O�w	C�I�\��Y�D���]�_��Za��A���g��Ox6��;q4擣W����Z\}�q�{^f��������C��\���FU��ـ�>[��!�x �F���&���0��V��(�]��I��7�*�x����\)��7v���GD�>N!��m���N(�5�R�_���8�5�G|j�C�x��k����!?�w��\bM�g����>u�lk�������B`�q�<�߃U��fwk~���<ÒZ�҆ X�`	׉H>���QE9�W�nٝ�R�7<�����u���ŗ�~=���,��^8���� ��w��g�+������������k�R������T|�X����<�/�K5*T��$n+��ҵy��
�<��Qʯ�����P��g�A��y�,izhH�����ߥ����<��"N�	�M6O^6yi��cb�թoQ��S,���M-�D�@&_�\QB�=�#n�x"�|�-O1�.3�ҫ!}���寫�(w0������'�T7��?��qw~�7��yy�m6�����l�֜�3%�绯BQ�����_&�q��9�O��`F���O�yk���~�n���^�֥��h�ˏ��E���A�B��7��kS{�Ò;�M�⑽?Szfw�{_��QK��voT�KGF�&����>��LU�ea�V���p�B�q�k�ڀ����2H�+Q�L���c�S:�P����_�$7���O�s��[����������������1���g�����wx;�Ko�i��D�itC�rꧽveI����{]���8[�t��q��wX�]c�\�%X��C|&,��VقƱ��q�U;�ٶX�J�U�=��i���.A�ϧ ������
��.j����ܤT�ڗ�[[ޙM\]y8ۮ��`v�]�ڦ�А�F��3~���8kD�:_���ɆЧ\?����;�*�beH9l�\�����6_=�|<~�ǭ[��MΆ���������2�$��l�z����5.%S�^|�_��c��9���#A���}���T}���5@� b���K�{�%ۏ�l�/T�-�G�5�L���4�����Rt�z\93���u�iz,��\h���M�Ie��C4\�)�򇋖S�ef�j��a��p!��L�L��L�o��йs��ᙇ��plI�@�͗3I�Hܛ�~��s$&�N�ߕr{�)�r5��Zb������*V�b����}"jA������﹞�h��ƕpO1kЫ�3� �#��ɹ��re=�!W�$O���:�3�v�xE��b�Ch��C��#�>�
J||!����Y
3E��gE�d�����x5�f�q�,�����3ĺι�c�\�-Ŕ��l��y����j��f�1,���y�Č���L��L�Z�7N�Aɝ N�����GTdt뗾I%�,gm���)�7Mf y��ܒB��KF��%p i�\���-,�x���-�����y�3��@���Ot��䌀�i�Hsm��7λ߃�v��ل�,	��7���"U:+�Xhvʈ�?ṗ�Uտ�����E��$��4s���_��Y:��7͆,�D:�9��6��]9���D3x$��[gUVBL}F:��<6��璯�������pK���Y~���E��s����4<bcA�܂���p
x�>���Lk�H�1�Y�I��[�mp`t�`��$�����M�M��Ֆi��<��e��ă�̛O�j1�J�#�ō[VK�"�&���Z���/
�
S��S($
����6�w" �*L���H�`࿷f
 i��NO�mi�0,軿/�ͭ`C�������o&̦<$�e�	�^"����o����7I�@��c����W��;<�������W�����.�e��L`jEN�=���қ-��~�ҹ��Jݖ*��"D��8?25�&Z�C��g}�ː�����?|ʳ��-�$����7'��ΦL���'���Y~**zJ�����, I�;��""�>,dl�ehu|�WHx+Q+�v���&ZTP`9{	�i4僦ܓ�.�<��N�"��Y�3%`)���h�y:4H2�̰��Q���=�Cs����7G��́���R9�͉���ʥ���6�O�S��1�l��d᭥<!�Ok�e,x�Q����}[���0g��m�k�%.o��?��z^k���:��ϻZ��핹�P�g�_&��p.���	F�|��Fqaǳ{&O���eX�z7�20��@�\B����߱,��H�܊֑��>eV�J��rdds�A��cSJ��Vȇ��ڹ�'��}nD���o���7C�{���Ɂ)M@� ��]̍Y\��<r�j)J�-P��5km8Q�|�>+����;�Zu"=�S��#w@��!�im^2�"�������� ����DǨ�&c�Up�줍����T����"�< �5�u��m�K���7�9#N�е���y�����U�މ����>�@����jH��H+�v����"6��nM�#U�6�r%[�iP���=� ����?��?ӥ��q�^owt���h^w�a^�=�/N��P���"�sjz���y�9΢��g��e�j���U�w`M�C�oƥ��z����I=^���Y����64\^v�sʖd�<�����\/�H�o|������?� m ay�a���υ����c������G�������D�͚CE@	�zֶ��]Q!SĲ+c,��b��o���ו8Xz-�9r}�ֲ��}�}����.C�q����z�g2؈3���yH��l�&�g5�m>9�D
�yG��Nk�S�2�mn�i����.��͒~&:��Zҽj�m�h:�$�\��B;.���B���me�����f�o�+%ռ�/b��:Cr)�JB�����j,�*@'�v
�.�;��a|tm����т�P�l��3�� ���r��81��0���u��k����*�6&��e����+Ÿm
5]{I˞�U���jW�,���<0��D5���X��-R��v<+�<��G�G�)լ�����i��:J��p��0�ļ����������j�Nw����q]��K!#i�X�c�_p���V�2��|�;������|�.�-|�u�=%hpt� ���C��ݐL�ŕ�7&%��r��,���l������C�|KY(h������ntV�Yʱ�vqW�0�uE��{��.��E�5�nr���O�j/l[@��'����|]��m��DD���z�c������XL�|���`$��o����+��}�A"B�hm:�k>�{M����ڦ:����=}��i2	��K�Q��d��2#�Y�0�9��.�U1F����7������`�q�A"&��x�kb�:�=��T�'(�	�ƀ<1Y>�؉�R��~��}���zqw��cO�׵�/V�E�ꇠI��dr1�<𧺯q�1�� �g2�J���x�sW�y(���g7*����w_�m��]��e֛���� ^����M�\��c,�6yf�X<p�λV�����Rb��n���ʢ$�[Ye� �x�w��	:U�s���3J��#��%d]3s�\�M뭭ؤ�|�|��M-���A��Z?��~�O���LP)7��i�]��my$�[}̛E��������o�����U�OV�Er��bٮ�erqV�6����/Y�J?��g�p���-o��)�'ڎ����޷S���66X�.�XU�i�<��74��8|d��[y0Ԉ�� �*�����i�ժۜ��:������$t>p���0��~�ߥ_�����q���`���z�q������G價�Ɛ���_�m�V�@n�:�8��D��F�C(A��a��@�d��!~���F?gi"F��,Z�r���{n���#U������ۥ��ۡ����P��D�w��	6j��L���G���/ʼ9L���>̪�m����7A��Q��G"��G�qb�R�٨�[��E�\NIh&���A2]xx�;k�H�Zo�����GN�*����G8'��N&Y�D�08��t��BNT2y�+�xv��h�53���QF�WVy 3��'+ڴeOq�^�ˌ�MS:HL=���$>�͕c�Ѻ{��[o=Jh����tS��6@=���P`�p���hߟ⧟��} ��e�Wq��F���͆Y��o�X�C�W-���}6�^]�#~mɻ���``�CD�!��Wjv�K~�ej�i����TiF�1+2�ÀUL��ѹq�j,Ft�F��ڽLr���
�q�s��3K[����T���O Ij4�}ߧ�%��Jq�^ڒk�$��kС\���L2�/5�:�j�z���(����>��i
��WܠK�WA� Ÿ�,�Y2�z�Y�r��.=ot�Gx���Vb��d �q� ������Rث�˰�G���[�8��ƖV���A���]Y��O0­�"B��+f�W�hsgN���q��{v���1FA�h����}�I�RQ�0���E/��&G|�?vk�����!�1}�hv�7�M�My	�f��Q ��}��4��,i
3e{�M�ryD�������P$s�Zr�Aѥf��4�����ܛǺx�M�Y�D�t;��\n���
Pg���%�%�řK5]|3�+��D`�>��*�W�nzbat�`����~���'�n��T�o�[�̍�^ל�u��:r"��א�Q��_�nلx������'A�y�AI�r��N���fZ���1�l������}����链g�f���f�̵^�^a"�|�za~��mn��i�������H��婷��X2�;"ř����z��P۝���
���~|ݭJ��Z1�ߧ_�_��xYm� o4_�p�Aͩ�3���9/1�r*�_��r7;��׆U�Wd�y�>�9o׃y�Cy��r�<�9���r�ą���N:%��㑅�e��^�*����՘�j������� ��"��˷�kB�X;� "�H_�\��up�︑YG7H�}ǖ��=(e���_��
MZ��R
�˴uBܴ�}�^�A�n&hJgM:�F�֬��;���.�.5��M�YC��W�Y���AZZ���$ѳ��אU{�O��>~�v�XƁ��U��A�d��,�}��a��˞�H�O�%y�ɗ��##�:���uũzO��s4R��؍m�V\x\��nMFZ5,C$�=���м��FQGŎ�3�C��~�T�/<Iw2�k#����� �2������6Fl{��@��>h-np��tݼ6�����8�c��b�B�N�_Џ�E*ȹ]|����u�4R����\n��U/���pa|P�!=� ����[UJ]��Z������Ƚk�'�
��n"'����	��k�QKֲL�����'#7����P��}�o<���%�=<'7�T���$�zK�����ɐ��h�S��h�2hs������_��<��#�v�j�9��37��ܗ�|T;��5l�#�7L	T���l"�Ȱ
«J7�:wk4�v�]�R�G��4�f�;�=��;���t��y5p�ΌI�ߐ�6I��C�	���ظ�ْ����\�e"�eNGp��b��M4�9��޸���/��-u��-b��U�\J�~#���[X���gݼ%�|s4)^u�x����<���;�֩� [d�9F���kj����Ca�-��&8ǐ�ڪ�)����em=��h=���c�C]'Y:��}E{�ܱ��}��A`1'���Y̱�:��$<Ƿ�D���n��ߞ����������|Fօ�Uw�D�B��˗�3-��D���9��<�|>w%ϠT���x��e)*�P����g���܌�-��)3�������B��/S��Ci�H���p[4m��~h�7�A�Pc�[��h�Ni��%I1,�ɤ8-*Z�N��28ˢ`��Ȼ<swi�!���r��R>k�@�3�!P�S�#Ҳ��X=�����Ij<#�\D��|�c�~��q`g�q�Ŝb��ߺ��U��a��K t�+��L &K1��29������{B��}ɂ�s�8�p/*�(�X�Жm�j�No�1�1i����QS��Z0.ٺԱ@�ᖶn~ݾ	x��`kǱkg}�faR.S����.��*�D�By3ο����E��E�)�|�Iw`~y���S�B��d;�`�0M]M���`�*t�Ŷ+�'X��X������"2��G��.��-?��
VB|�=��+S΋�Wpa~�'2��A2c�5G����%��PU�@^��wE��G��|��3X�j�أ���ۦ���]��Ph��TD�wơ���6�������Ec`~Vj�� �"��n�er��۝N�M:Z�4���E�!��,�r1F�KP��%�I'�|}��:����י�{lR��>#������ź�wg͝3�^3�Q�5�:$�]t�ֿ#��73˵͉�}
jݺ�@r�����ߦcĆ�"�\�[�<���岲T���.IZ}���#@Ĕ>���志.V�7�^l�uk�G[7F��!�;�7�d"=E|����VG*�>R�h��������ψ�w��z�����*rD�W�Ȩ.MuT��I�0~����� lؠuc��@%����"��%���S��'� �;�wR���0��L`�O�a�<�ɛ����_,�$�}�'��A ���z�
 d��4ZEZ�������8,���R��*=<9!�\�)�[�Yg
�#�ޫ x�?��qY�'����t��PJK R����bjK �0�*e���V�+��g�L�`�Hp�ok���HYkv?�	#��a6�[�"�3�I+�oXi��=v��۵{��6�C�X�WF>­�O��6�Leo��+�ƋI����{g�Ư?YY�u���x����O����B�O��H��_>�8|4����Td<���f���ʁ���Ȼ�B������u��2j�^��^g�c��X�"Q���p�?���:��)��n�,�tl�vc��)�����c̟��[��[H��+';=�>!����c�H����y�m�[3e��]�I�;��,x$����\�8��q8��W�w����{f��O0�r�O��pH ����,-�r)*,C_��D�8��a�a��Ѥ���w[9��7E��~ ��)��J��nT��l�6B��c�'=,�D�*����
� Ʒz���Q����W�
|<Ҹk�w��p=��3��oːƒ*��ץ�h~����5�4y��U0��<�
��\�L��g�߮�>Oe��j�k������`I��KN��*��fL�k����=� �_	��.�oj?�� r���"�~��|ǓȯG�!m^��J	��l��"_�9,�L�<:�)�m���[M�!�Dd	>�����N�k��ߺa󾐩k�����Ԧ�>F8�����S��ŋw�6���b+�p�DC���o`h��͓i��Ҝbd��?����ڇ�=='K
�����.|���*[I��!<�S�"+���ɦ4���r�`�p��s��=���z��?� iY���t�Dw{wYp/º=�O���:n����A�N.66�PUy��j�g�H���	���70)�ؗv����$��5�w �����..`L,�$[��]6�oÑv&��EAD��pVY��-��1�o��"&/��đ���A�xQ9�>�%��n9=3��\m�ݷj��_�{IT��/�|���Rw.�����&&��k].��5.7$oC���ǇJV]^%K���|�@u����6�>� �4�s��+�y`��K���c�G�Li9�FgXg�`��g�;UJ�{�8J�=:��Uj�dOX��"��L,�W�Fe�p�Ǯ�����.D����O�D} ¤&�5"#<�%/���g��6����������tl�G*���M��*y�i���8���5�D8X�Fc6�_)�'~�Y�L�ل(y7��"���S��<���@&l�m�
M��r���Yl�;d?��F�����/L�.S��� �T�g�;�$��wX��o���O�w��[/!�u�� �������/����Ut㠭:5RP6D>;�k<NUH�Jł�|�$ZiY��T|1�-,�WR��vܧ��Za��
Z<�����[�c�����{Z���~(����-��k�*���2�_��̌Eч����O9X�o��@�v~��5Z0�J�o|�I%7����'J�#�b-�_�֋븑(����2x�W_�<'���$�t�ZU����]r.[�]���?�Y=��[W��>�8r���Dׯ����g�I�.�H.�!zPAx��,�K��aO��T���x�&Z���MO�� ��4�k�Q�g���2��/rv_�No�3�
2�܊�]���n�ֆ*�+m�`0^MSm���o͸>ݤ9yP�/�����
.��Y�$��/�2�f��a�qZ%y�5Yd�m������2�%m!�A���K2��x����CA�s�����������'U�l<���k)>�NM��[�5�U�a��y�:�[(\I4���1Ћ%���l[�4a��;�Xn���
�:V�z\�,R>��D��P<U;�,I��A�9������i��y�=t�G;�-�&1+���;���2��
������=}���+�lh������R6��Ƴ�|y��ދ��jin{�*�-�:\�P���Pnv�3����;�%�m�f���k�\&��*�P0�9��7�(;� ��x�*�,���Jd�5�߰�N�=~�Ok^�����@]�'���C��w�;}.�ͥg�/a2�zN��{搘���e��б$�����N9�~:`����n�q��͘�{�^�ɥ��aRR�N��i�:VM���He�=tzA��V�ȫ�.�)nL�?���Ù��b$�L����m mY����+�(R�}W��ʛ���*`J6cn�--$O	���~�oW�~��e㦧a��ՓJ9�a��e���!�%�y|"�5L	�^���+CO#�$o�����\�Qw� �	�*D����䶜�{Sd^�;��70
���{9�p���܍i��$^�\J.�74��Y��n�Cb鸭D��3JC��Y��9�0Bh��&�����2&��m��ևY�������
���B�(��K����������'
���V��wI$��<�����T'�����\�*1�������_vRM R�vRLkD�:q�S7��h2	t�}� �G�D�?3�U��f(�0��-Q��e�!x��y�.��y\��ZX
^4�2�o�4��������\�1�=�s�pg@|{�������Th�	�r��(,mJl9��f��%)t�ߛK�K�n
�c_'��zE�
#�Ŵ���=V{X�~(6/)�F�de�fk>��}5�{J;!������O��f�V-�XN�D,b�C`53r_LW�c1x����dk~�as!�[���%r��{�� ��&x�Z���z*'/$ُ;++�p��Hf�x�p\1K��7)�Ω��U���{�|_��i������E�����ɺ�����M^W`�N��>�re`c
9�h�'�ANM�Jn��+�a!��7�G��J�^��^r�3A���ه���=`!�gy��	t��˔X�v�5����O]<�=��u3��?4"I��+� ��,������:q/�0r"���L��\2ӆ����~�瑝x�����X�����!K��Ӓ�.:,�MI�Ij`���\�~�e��e���|���
�����M�SVF����~=��̧ΐ��&� fv9�t���r�,?�hdޡ��h�n���b�۬I��Ÿ䬔8�����rAP�~��;�aʼ���&�YXQ������k�H6ex9֏{gk��W|x�V�01�U�/��)2O�/r�ر��Τ	7eX2�m��z��S/�K�$��S�X��$�q��P�}Ε�x�q�A��m�/�s��d���=Y7X��q������ӼBil�>��LK�J��G U~\<����Ih�,�&���q)�M�uu�M,�&��]j�-:Ԭ��6H5�9<l����wS�D�H����7����j�R�����6_P��*g'c����`l[s���'�M�����l��Tz�\Q�s���H�6���B2+�Ɵ�?�#q���Ï�R�Y6�4�����}s%��SèڑٛHg�����-Fߦe�#�G��R_q�A��ʔc��Ј��k�LsF�MqY�� �*:^\��|�Q����e�x���O�$�(J	9��3�h��5�2���<"oҩ&���~��t�+O�T]���0"�a�;�*1�R�ٿR�r��r��G����P{P$�N�T�����|u4����߱[�ر,_ӵ?/_c�|uҀX��1Z��3�:��byՌv�i�%#������P�N������&�"�/bk��ah��qGi�B���G��[���P����LJ������)��@���ͲP�_ǝ	�ePHL����GU��I���s�����b��8�[w�r� ;F�<���'��������<^��?��3���%#�Ht=bk��b��.�
P�˷�x����OF7�rN=�����w��"ǛX����W��!2upd�dk7�?Z#�~ï�@�{?�e�"��8��Q`s	���ʝ��b~v�A֔�,g�f����B;��c���T�&W ��ߪ�(�^3��M�97;?*hmU��.n�[��	���h�߆�B��O�e�����|��D��	�^�qJ���\<�⟫�m����ױ�қ�2K_׼[3��I���_�&{	,SY@�n�K��g� �.��,���u@Q�wwA.������}`�Q�ݔr����˓�m�Q;�LN���9~����� ��vl��GD�@S���C�زK����G�\n{�� Ʊ��T\�I�-���˓m,|�7�Sm0�%�F�К�!𸜝�����T�d��%���-A�B��2�O�j�/�M�ϔ�,���c�[Q��7QmV�����o�Զ.� ��$�w��݆���X�G"4)ǟq�R�c��Qy|	U����j6X��Wk��͙1N�r�H�,�4��D�R�[n�{��B�r��<ZH���|��2 _o}�����%=wS~;*�����rYpZ�b�)�4�$�p3��<�:&�{O�D�A�vڟ�_a]�����`���_"=	���oϒ3�Ź�-f i�O����!�Do�H#4��%���:�� ���E�u.��ۣ7`�b��zJ���,=9!:C5�n�c/Zg�/��G�,[gF?�~֧#��(�"c�����[1y0B�F�-���Nb��=��Hɨ9e�&���w%A�v)�1YC{>�,�x;��L����G%��F{4��-/r���������C�b��������5nȜ���NY5���0����Ty'�٨��Ui*ϱ�%{�S
��n?i`$�:�y/������cdjgfE���HڟW�Z�� ��%�K6ZA��d�0M�y�ar����$�pV�Lö��.Ϸ�J�rW�({ȥ
W{��i*�{����eB���㹿�V=�m��}8��xw-p�>�`� .<�*�
ڭ�6;T|n�O�� ,�i
����C���_���3��ೊ��،���Q.H����F�=2�䏞��J��+R˿@�-%1\�Br1p�K��K��?r�/"�D��/O�8� p�K'R�x����!�HP}�ߕ�~�o?�z{��r��k(4�$/�d3��R�7N_u�d׮�n�<?�|:+m��6 �7�2���v�%��+���J��M%�;�$4�_:�r'�����EL�9	-�����˄��]jsa�{d"&���:Y 
!64�*�#��B�%UF�p5�2���M��~K������цkC�/
���#fC+�
"�(���Q5KRm��3�?J*
�
%��و��RD]�rd�+&�`H
I}�hɎ�#6�$/I�N�]>�om!O=�µ*�/y�p
���c������+�]`�'�nF��¥GF�k R66��jF�)$���"$8���X�M��=X�@,�B[���u8/�$��%�^9��Jj	 >Y�>��|�*���2��+��QywzY���ډ��'M(��Cԭd��)�cԢ�J.�jk��Ѧw�C��l3�ua�&}�	q��o\�J��:z�U�ը��|+F��&�0��OT>�\��*��m^A���En@���&����`�|�df��:'r����nB��ҭt�ۗ�������	�1����j��?������U�,�<1���]_O������G��$����{��>��0S7aܵ���z!�����Ok:�����/��7L1�]X;s�����'�C*t��.��f�x*z�Q�F�$���ϲ湫����W�9�'���R��0�ï�
s�#����s���p��˻%y���;M�`ԟ�$�w��n���zS[�&�Sf�.Ā渨��*�z���ts�ޒ��O�����BI&n���^5hq�x#�J�{i�
�T����Ģ��0b��B _W���էaW�S����i)���Pb���
U��+V.��\G	���ܭIOS0�V���TR2��:D�R���A ׮�u�v�rާ�QH�e6�K藠P�飯����7�M��d^e���ۼ����cxp��w�����Z�b\�o����
P����L�\Ee�ް�_���o�<Rs���&��G�E.}׌���V彴p͗��k�P�nˑx�&?��нo���lQ�Kj6aGO��i��q�,m$�^��\9>*)YYd �?牪Y3{%Z���̐��ꆳ���]r:���@�v��w���x��Q9jC��
�ۖ3\٦r풖m��3��jT-��G���t/78p���׽��X'���ͺ�_���ͫ�^ײs��zC?ĭ��]�@�)Xf�d�����s��!һ�%�8
TU�@�<�v]���7�[���-�.,>w3��`d�����6G<��k
�-��e�䲦�8���EP�O�-���"�`��ײ��H���ן�,�&��v �N�)�m4�ff��ߧ��Z�d{D�7l��s2�1
�k���e}y��X�>"��X�>rs�6�X�	`R�+%㐻V,��`�u�ʻ�mg�PJ�MX�1�5���Pn-�u����Ό�{زYȭb��3J���*������(̀�TO��1�O�/�3bi���9z-����yv�S���*�{��̖��e#���b���-����b�X���/p]���H-�/^� S�16���m�]d���ޓ��H�v
�L	��N_����6ټ��	\��Kh/���z����bqz;��c{U�\T�﵊m;9$)1V��(��w��M\z�/����-��gq��Z.dό���@��vU�L�*����I7�8��� ��p�o��07�1�(]�FQ��P8��= G����.�Mi{��e��� ���{��]��+���x�6B9������em��~I�@��{��%��r���$=RVꖖ}r�.���q�=����+d�;���ֲ�!S�]�>���y�㳂V�r��]��P6��'d�L`�4~���6�g�Vs�í���:{]\��g�,'Т�;���ʇh@Eߘ�9Z<�&��JU�qT�\E*7!`�S>�{Ȣ#�5�@����w���9J��N7��Ed��L���i����P�/9��:XG�	�N�g�s���=�1&���A���H��+�Y��%[�a{�A`�E2x#�d�p���bj�o���W�4�b���˝��H�,?��v״٤ڮFż�t�k�V6�KN�p�����y�6���'Dત<����M t�cѓh;$R�z���2���+�Z�aH�Ҝ�_�V�遘�تt_Xw�4.�th���Z�\��I�uS�ʃ00m>^N�[j������D&�G�ف���]���6f3�؞����[x��ɧ*��{�o�g	��Ѽw9m~��Ц+;�D���(��D���S��|�:�\o���������KN���ҙvf_	�5�"�||�xXЫV�Os�
��$7']�<w'��1�H�+�IIz�ve�y>����S��X(�1�Siw{#�����)���C��6��eU��t���
����c�%3۲P<��T��qAr�J�k��gd�|nE;8�:��㽗R�Ue�J񭀈n�e)1,�=�[�gz4d�AlI���7i@�Ǡ���5�|�|[Q��Q�v����?p�b7O�L�U~����*��P��ÜlA��I"�VHrG�
 G$�B	�` �!����f�8��1�,:��_�+��>�	n;щ{ȇk��8��A�����!Jbr%�e��{0�����F��2D2��1�8�Ni1Ü��VW��[25��Dg?��;E��;�*@��Z4�
O�n������Z7�Q-fg3/��ɶ��J���ul	�&AM�b�n��v�X�~��T)1PCS��+�ڋ�1Q.�/�c�����9+�v��:���_@�Q�7w�R�'�ީ;z$��pT���P���~��H���7|�H�>�tLO���`�=��]�B׼�r�ˤ���G��]�C�a��Ė@H�&�u�Ot@-�.�\L�P�QbP�V�B/,����������6r�"*?Lԍ���*���%���Ȭ�k&c �C���R�z�~�i�~Xƌ�7?h^ݱ��iasL~�/�o-�G*m�w�������ќx�,�"���o��r�A�y�ߘ��u-����o�\.>T
���Xs/�?�텔�t��I!�Q���!V�k�����G4^�^��]IfЦ�#��4�ڢg_�q!�]n���_�~�� 6*�'�L�Ɓ_wfr�*.���
� �ݧ(�LIscۅ�$����*r�F�N�38-2��:i��E��U���+�q���[���Ȧ�q��yK@_ߔt����Dd@Q_t@�>n�(�![�0R>޿?Fz���V��85�X�K��V2;:w )�X�����d�a5ٷ��L����v�|�~��>�2�P��pc?�R7��7�c��@xW�&#ݶ���丟��JQ���\����A0�/��d��S��B�x��m]W��J�b��t�5v��8�Z��uI-�;�#a�c��<ٷ�ɀ*)��D5�$Ԛ:{ �؈:~�$�D�d2�3o�����-��چ��}!�OB_M�Gk�+Z���,����
x]X%#	2?�r�U!��_+�}1�&_{�E������t�P�RGF���2��i��o���NΦ5
���x�����5��ə���I�k�ez�r�og�6��w�3vxT��ǰj&�]'�����&����P�$g*�����8Z%�XRX����ސ��5��QS �7���l�7�n�J����ʜ �@�	�_�;hU��3� ��&��Ա��O����B����V��k}��>�0I慚(��Ч�e��/��=	q>>����Q�k֞�r�x�$���������I<�'�CO ���;���\�a�ɦ'Yt$���C�@��D��+�#�3�c3������2]2�]/����.%P�n�Xtl��K�������H��\�E��'m뽡��d��QR �Q�m�C	&�xT�(�/�9�74�5԰T1&��5k�8}/w�\s	���\D���9c|��� ������o$����S�	f�O��G{��v�dMXgҾx���G�2��D��<�7�
u��n��'V�U՗�5 ����]������꜕��gǶ���^1�{9Ĉ���=�3;1� ��ؘ��N��FT9;�*D���WbƐB{�q�M�u�i��pՂO�1�O�n�3ڼLrC#GN�W���� ��s|ԗ�4?��t�4��4�i��_��߰/wd�A��q�|>ye��'è:��U�:���%ٛj���/�o5r�x�h�\��EH�=�O�!�m�/���H����@���X\X2�KE`�.��S���:O�

��|ȝONnA9����w�7a�q*������|����PMm[�T)JQ@����� �I-TE�-�nCA��&��PC�K�%�J@Zh�?x�����{g�19��ךkι��|���R(ԑ��WL�8��Rr4��yi{��l��a}��Sc]�I /����$��栮<��{���Y�oLs�:��k��p�m�����A�V�.�^^j�e|u{Zފ8����Z���ʳ�����3�dh 껼��^'K
�\���?C�FM�����۷m�z�Dބe=w�P���:U*��8jqR������j������Nԝ��?GZ�Y`*���.��_ʡ��%�ی���xJݾ8�2�������E��s7$������.�S�w�vv��h�o��f,���4�F�If �^�47t����ӓ}�a@1���7�hE�ܩx�<D����cT��ˊ��F蒜A�H��4����g֗�q?��Vt���ۉ((�t���3<J�5�T�Ay���+�WD���i��W��������/�)%��E�I���^������o�7��B������W�qG�#
Fx|h��[�l�ʠN�`��W����:]z�ynJ3钽�	Ѡ��.�oߤ�g����2�^��"���"j~�b��Jd$�.U'�>�2�u���vv���?��(f1��
g�?q���C�CK����]B@v��0H��BD�\y��x�^��jc�5�%<�� ����J�H F7N@��ۿ��>��㐯E�Fo���{,j�����课�O������,� $��t�8>xq������R��C�G�����}�5��ž��I׿�S\f��1%X���p�Rp���me�'>�&�|��(�����h�{*c�Y~pO��JK�w{��(��c�TlFi�YS�	�ˆ
�F�fM��u�)z���{FG^���[M���l4b����+�6��C8���J�Ji�I�e��jg]����K|ictku�h��^�_��ʙh
:0<�HQ�J+q-�		��� ��R�b3�i���-m@&uyi���W�C?�=�=T����,�
whxp�DDX\��*�mjQ�d�����HՍ�F�$Q��������z��G_dvP ��q~~���@|ŝ&��U���.8`$j�xNb����_����gҐ�پ���YH�_֔��C7��KE��S���J1���������g�C��|Oʚ��{�˓�P7����Y/+4�k2R���p�v�P�wU(Ų�R�q�ypMgw�	N����i���m�9̹o��_+���Z#ך^!���5��1x�̹z:>^�����	����ǯLTD��Y�Gv�nNP���G1��+x������Sv�>�Vn`%Z�"T66�G���t\�	���E��K����p���J%�?Ow����o�k�1��BIs���|�g�"�.	��k>�s��>=���|��h��u���T�>u%��8a>�m��$Gy��o�oi�����g]����ק�	���S��9E7�݊ "�D�+���hi~��/����������١����?���m��gx5
@�Bڛ���.�B&��&ץ��~c��d.y����,Ä�߽��{1�}�K0����a�B��1�\���ڳ�4���.{}�>��#��a1M���v�N��s>��%���:W�Q�1��O�䞋���VM�9X����n ᛴ�f�)yC}r���i�O�),���g%�A%�Ɉ�*9�We��Z�is���y���\�O%����=��Q(�g�9�r2�9�?~�n(�R�%7�����B:G y�z�v{L��ˇ��<��I�u�-�&�z+��������ײ��_y���E{gF��Z����9k�7m�eU]�ؿ-6����\~߷5��Ha���'x��`�����̇��>2��_�
���t��&��Cn�,;��Ǥl�g����O��ƨ3��[8.Y$�<&����7������Y�%�:�������Ȏ�?Q�ɷ�٥�����*6f��޷�(��i�ﺗJ�$K2�ܙ�r��U�o/E�*^�i�|/<"ޛ�3��C3l/�Ft�Y�Jo�L�>�`���_+ y�Y���g��h�%$��Z��3M�щw��$_P{� |��#�4����}J�|~��ȥ*[P&������4��_%)��Y�:�Ȭ�C�0G.x�Z,x�Mx���ͼ�+�G��dR��K�({j�G��C�g�ʛ1����@-��� k����T��+OB�>���̷x�d���eVj�j��ky��s�<��vi��y�E5���+�%t9��(K���_J ~q{�~�2%�d�K� uׄ;gS"����
xd&��&�pzsT]�Oڪ"�zug���6$~$�"W�?�թ��ȏ�u=�{L*\�N��?w��s���^��g6� ��d�!���7f8[�;"��}5<�6�o�E7a|���9�zԣ��5�OlZ9�q��fz�(u��Um?�x����i}��f��ßW�2Es?!N�D{���^ɴuq���!��a�s����}Tl��vb���Kf����<�W*���	��~�@�Fʶ���54��*!��Zu��w���xxޢ����ᭋ�1Y`g�;a�R3��	�i	G�52&�����<yb4�!@ĖCW/�����d��Q!Sm%�!��g[�����������{*�Lg���ĸ��K�<�}v�c2xHF}p!�z����#�Qx���R)p��!/U3�|}��3��f���i��;�����~r�hEĳ�Z���U[�3}����2u��d���e�Ҭ#��9*���3�Y�*������Ωf�&��/�_)���E��8q�����͛��1q��L��2�ΐ����s�<���!����>�M�T��?���'g�Cm�q��������Y�{��я������+e�.�1��E��W?���L�Em+���si>T��kW�Y�$ ڣF�`�o����U�=���l�+޾G�g��R=��k	��J1�3v�kd�J�v4<�Aě��QpJ����Q	ٝ����9�����Cye�/����gϤ��PT���֓ݝL��l�aK5���V���߂�T�T�|j�����0��|E>�Z͡w.'e�}��|_C�Լ��Ϧ�&����$�a$��T���E�<�_��צ�𓶨p$��u��t���<�_�k% �!S#za�<n͓Σ;6�Vm`�bڹL$��U����g�g�{/-�W�:��ۊT�S.n]�6�wn��+��F��i�;��(Y?�.��u�\߸Bz����=�DanU�
�v�-���M�R��Y�V!;������|��g�aUy�иKS�x��wvtjN�k�"��6L]�X�<�O.ʽrC�7�� �J� �o$�\��p�$ۂ��1�������x�,]g����t呣������/��۽��ۉ�\�kN���sw���,[��j���2�ܥT����.�R�d�;oWK�MR��~����x�6&��֔�_���7����Z���#��c���7��H93oo[a7�����P���L�uEi����PO%^����h+�q��<�L"zά}g��%D����3w���HҤ��9�L�Ui���țb.�Ԇ&�T����P�l���U{GG̱x�)��9��s̪�5�S�\�5̐�5��/Q�{ϐ�Na�kiH����=+U��:�O�4�n����>&R,iW��(�mhl�6Ԕ&�5���?gC�ۼȦ\x�l4�l3f�%�#֭����Hl3z�����4.>w#��߇Y�ntQ\
%��ĐJ�N�����v�E�!��[�[Bh����Y��a�-��W��WR���d���	�}_���zW���W7�XW ��:�J�Lr~T��m��oҳ�l5G54k|�ƹ�s�6���H��I�]!������-���1�0w�ڽ0�Ai���B��F�G�4=>NW���?wy�j�Gv�uă�sӗ�E�m���~�`I�����[�u�[L�ݘ+��
������<�BzB�i�U��[�@bq��5~�{�G)l�"/�,���y_��̹�Hv_�YhVZ����&ĮO^Q��c��������L3�rx�%��5�,��[�a��c�6Y�g�4���i�7/�y���z�dVf��5���mM9]%�l-P�v1�f�aae
����F�Ñ���-:����1N�����b�/;�߻5m}$-ݘ'��1y>h���L��{���8���4;}�$�ʹ�~ ��#2�dia	 �V�Ot�{�_�b������H�Gk=�g�LùE_,�h7��0�Z�_�x(����3�*#`=��q�S�g�q_�s�'�~��N5���0v7U8)�t��ٓ��9�����<�y�ȳ��x��!��xoX�յ@����.�&����yb�mO����pXu�6џ��9�y�u�7���B�-�<{ߑCM*����N��O���S��L�Y�4&�P����ֹ_�BZ���?nF+�M瞎�mp��V�����n��tL<g��|O_Vv���%���]o�8�p��p��21z7�i/�k{�Z|Y��W~d�,0?�t��'WH�����O�[ lb�iU���v�e8��_$���4����S��V�&��0X���gx�*uqt�A`���@����$��Z^~OA�ā��x���]5/@����K1�b�gz�k_��ήD���&_%����Ɇ(�=����������;\,(:l��@1�D\s�<or��۔>��L2����NcP|�^Jq[���7������2����.!lDm܆|e؟�XGz��#��u�!��A�N�ԗ���#~e�����fj���M.uq��̿+b�\O0rT�}*<韌����9��i��FP�?���0;���}lU���҇�%-/,at=�uNj=Tp���@e��@i��W=�<(�ߣΘ���㒷t:�c��%E�@�%�՟���L��(�g���Z�/C���|��5(�����Ru�x2�:�{��\lq���L'��˿�D����0i�8h�ER�UƵgc��?c�#��TM�{r�6�䬊�o��j}�,}�]�b��PJ�rw��N%L I�������?wy0Z�H[y���OZ;-'4"�(}I"��9�|�U�ك���jb�3�_=�ʛ�/9�>o�0�M��J������M�ț5���D�+k��b+��_�Tѥ�8�=��]����g���(��*����]��/��}y��d��7��%�q��bޜ�Rk��ɀ2�Jk��K [4��me����y6>6�O҇|L��]�nM��yH�-oWgi�(���b~���E��.���S��Qy�wʼ���o�?;W��0�>�n��v�zQ�?Ejw�pƢ�r�?(9�kVh�r�)��_�Q�s>�h߂7�%e�#�U#ܜ�5�Z�k~������V^��7���	���|�9$�,��7Մ	z�ԅM��Y�y)g%��8���Ն�P���� J�A@1�cW����CP@�Q�K����}ʂ�--LQ��U$�����/��	5���U"ǻI-(�Fvj$����*����s�F�ծIԳI����.�V:mʱʔ˾�+���x.Kt��vg�{5��N�"���A��5y'�;ט�:�����Fdz�����8p�ݗ�52c�h�z�G��
��4k~�_��Z�kX�h8�,xe�~��o���S ����F��F*[��L<�_�k�ְ>��J��W��k[F��j<��^`C�����6�@��~�K�҈��py�&uuPk��l��R���G ,Kn���?���[��1Sm4�*��m�Fׇa�r�ua<����WCZ��vj��6��Yi�3wҨ/�Z�<U!�63��% �?��;�~_���4�@X)ni�}f<R�H�2��`4���dgf"�!3��/OJ+��۝#���ܙu�H�Xt�c�"����Dz2�M�-�5+��+JYp���%Qh��x�pr��fJ�H��]0��x=��BN���<o0W���1�
��Q��H���)�?��\б��,�<	4�^�d�Q�����ɖ	:d�Y�Zg@���e����S�������*s'W�����C�G�,>���G^~�	�������5C��em�◪�����L��nGEk���G���Qʲ���ݾ�йc-;��,D�@��Y�x����~���iގA���B[Ŝy��x�8U��.B�/Q��A���}�h�c��"� �f�Cw}|7��/�f�h��`��a݈�I���j�Ș���H������u��3��6�Υ(��r��#���q��������%����k��j<��;�F;�S�Ǆ5�{�xL�lDH��9�2�Cڝ����q��	\���w�}g) y'���K��	���.�f$�+ݥ�ұ?8����ȏ�l��o�"�2����$T�^J͒7��E�kμ&'�>Ĥ�Uŝ�H���>͆u�y�
Oa/�v�ZZ��v�3�Q3���˂��t��+f�Ч+�M�;è�bV��j	���:������5��_��opOĞ���py!��oޠ��b��}�_���ύ�>�{��@�}��,����?�D��߮j::5l)�\/;�P�)+���ϫB�w"��~���~��N`+�D.T�K�I�_%E�w���/8��p����em:��g�T9��ϴAA�Arn�YH}ï��t�ic�3O�W���iL�����ޘ��Q����fh���Z��ʄ?�(`l�2,@�M�6-���p�zH���p��M�s�!}O(����'	\f'bK�+��pa�����)A�|���>��qעU�d��������]K/O�ۛ7(�����8�V-��S�FX�J9���o^ �u�J�A�ڲ�_��c/��`8\2���$aX	�gbb�=���9r�z���)��8�Zx4���Jo�L"����O�F\��K෋���>C�̨���3�V�xx���	�Īy�ʒ�qY@�$\wqyL_A����R��~`R��S3i�Mar�.G?�x���$�?'����(4"��ӧ������Y:�Ag܄ La�¯�2���؏�a�=�paG/>؆[��'�~~M&�,�j��_di.β^O���O�4�Ms�6Mq�CWY�$�e[� M��	�oG	� ���EԶ����8uy4�i���\'%�1꿐���ywÊ�=��c���S�OA��R��ok#n��o�ᄟ��h����Dgb��0���U��*�]�n����Λ=�P�5d�1"�g��"�X�w莆]wy�,��+k�����n�kd$v��c���5z�3��8;�^�E�B~,S_���ϋ3~��'S���zp�KV6vV��K�ޢ�xm̒�S%��1��^�������{���k�Up�PQKɣvͯE~��R�e�3�����6�w�l{a1���$��?I�"èD��?=�i�:��~T�=�h^|�׋-
��F<���1	��ܩ�MRe����s��}N��3����Qt��)�NO�B~Ѿ �%���D�"�[k#��~4�8�c��*S�^b��.�%����
��=�5��sk+��$���y��
[�p濗�����u���
�F
��D�;����������m�A�Ecid�-�>:3 9W�/�N52��'��/�R_S*��G>�������1���¿y?�[{����7�F��/$,�mO�kC&��G��tM*�gP�XPy��ˋ���d_�~1У��ȧ0��bw�JkO�����J�ee���VZb^t���h��Y��Q���7���K���v�z�𵮵�m� I�k����/��z'4f�"���L	��&ċ���$�WB¤�,�O�?_�]sa�a�z�Ɛ�>�i���-7��@'�~N�����N�hT�9�.���mĚ�Rڅ�c��J|r>��=����2|]�R�b��� �`�h\�
H �Fn��z̾M����gG�l����P;~=D���P(�W���dCQ#��������\>�������޺.������r`m�7���T����g��e��56&K���/>kE�ðA�u)m�Nub@��	ݘ�gG[\�eĳ�����"��L�������]{j�)�ms�[P�"tm*�[ $ָC�t�K�{�35�Z>3���`m�a���ɺy�����tG�߲Jn�[Ӻ(]`�bJ�1��?MF��n�+�`"H�8�}��34��tG[cX����G}�ؖ��z��@P!�R�A�:烱�/���˗����OLB�)9��6�?#��Y�N������o��5CT� �0�4����G�c�#�_��m�����~[D���B��]\ō���F���P��g���tR���sy%I�"v�$�Y��X��~0�k���1�m�˹{�5h�pԝ|E���CX�G+��6GNK�j�Y�j8g��xC�x�W�FH�B�O���忠��+��c榏���Wg�	��Q.����a��4A�}��"�B��C��C��{�IOU��x�ޅ%oU���R�w%�^��H�G�'�Ey�[�II�/A�X��S@5���&��[c'�a�_^!���za��gZN�6OƁ��9�-j�NG�v�	e�Jz7i~�/��&�x�/��V��Ba���K?qZ�U�7��79�����T�N��}PIӞi(YZ���E�Ԓ/s�'5��Y���l��L��|��&�:�<�Jx�o*�6�����v~T�j&ni_��&@է������-�}�TY���k}Z�����p+�!����� *V����f���75���m�5*�L�W�6	����O�����%�������Z�Ձj�?������=�c����jh�ԡU��Xq�5���U�9��|O�=�[�$���E�z�eq2�7�!w�����y�0e5�I`��݂��+������=Z�5C���=��{������C���q��
k��aB�m7��`�9�	n^-ν�'R��N{Z�`W�t4u�����p��bAj��%t���C�۵	��1�����SG�I.��GzJ7�<�#,�{`�7����Β󟛶K���=�{�k�$G�u�^
��Z����{o�8���'�2�z� mV/	G�0�d�Ȣ dU05�0�"tA�q�	�W�Ը�
�8�݉��x8�KR'��f���RJ�T/��9���R{6i���$�0)�,Sb1T��r�4���MV�����*� �7�R�9@�o�N�"��Nh�kuǀ�-?��o��:�PGDT`\����D�o��
T�|�>��.B[�̸(���₦2����Ad����׿/��F��n����ǀ�.�4=fJ�N �)����>��^���>	h`Cv_��#^����-�]��k���Q��N�Ͷ9��Z��|#�48;����^��2�ݘ#�,I,�`jR�~g����\���E���z�@Y�Q^����̿@D"�}F(к",-�Re���R!Մ�Žj��T,W��%D�\�+����7o`4FyX6��.d(�@��198�ꓨ�A�zL���[L �' '_@�|�f�"�jPG�I���p_��O��A���f�����3M�;���2����ݩ����J�a=�����q1��rW��`7�.M�(m�_�SR�|1ډQ_/�ZWL��Zzq�`Z�p�Oi�=�0v�1u��v�S������?�9��P�wAN�1�Cwa�}���n��.ѭ�gw�؎.<�J3�����'垨:=���>��p�)kE�����	+�a�)��ԳG�R�`[Y����e�j��:��5�r)�`��E��.�Ĭ��4۵.g'���Ύ.{�!�0��~������h��|w�0���[4���b�!I,� z����@�K��Hӿ�G�U�<���m[=���;�5��'ގUA%�$/lu�(a�G5P��k�N��N�w�K��'0@^0�������f������g�i9Ӫө�4TؐM,�W�.���)���/��~�;,�7���D/��/f��L����]��a��B�<Lۂ7N� �E��B���%���J�<����(O����p�k>0i$�ܫ������Ӆ� �G����Fk��J���Ρ�I֠�O�~K���V%���oZ]K���&��/p]�7��՗����	l��.�Y��N�<��û�=�Q�f��@�����񩡣�wы�p�Oo^|����@�j�Bm�P�JTyCJ�>�B�se�%�ĺ�Dc�k���t����+��43*U���v9��\{m5�iH^oo�cQB�����B���^���9s������q�nA�ԣ�F1�M�YP��pg^h��&������|�Y#]�g>�����ط.��ؗx#L��觲��6���X���{��JSXv����{��
�𪇪p�XM�L��n��5{p㧞��֎��<�BQ3��"��F�}J�p���U�>P*v9���n�<���yD�ը��~�ZW��9p�fˣ�h��GC'�X,��X2+�8-�N	����|%�c�����UG�����B�KՀm���p3nA�5��vY����
�
��;��G���w��^����:tC�T���f�vIO���S+SJ_r�;cq��Ό�����k�����SW�3pF�CƼCY�*5	#Yv����OQ�	5�=1G�kE�7e��#+z�^>����aߟ\��e�r���j����[��{�+���[B�;�7��I�@dk/ͤ@C�S�u1�O�����9���Ϯ��y��i�H�Hǈ^b���$�P9T~*�&GK��O|��O��ݮ>Z-�="��u�X ���4��9�����ݼ=��)eQ�>o�rzx�@X�/6-80��5<*=�j���|v��K�uc�!�46E�;�*FA(>�U:�%�"�r��O��CRA��y�aw��X"WH�I`P:�Fm��|��0~�l>�/U�SV�������	5�^�F��Y�cդ�DOdr�*p¤m��<�e
0���rH���Z���ĝU�MMnuRM]5Ս��IS.�c�i,���{sw�]/����g*jJ�H���ի}�K]�����bFL�����j�S{��W��x�T���lJ5v@4i.�~@k�g��&��/�?�j&����*]��:Vk�-.4�ϙt�F�Vp�z8TO=�޵��zJ?��s���`�� �7��-�TV�~N����%����-�
��%�+<����c	2]D��hR(��P��2!�*�eܺ��K�#O�[-�g��A�|Bh.�l��rއ�:b%�Y<��UU��BFC��c�
���尺&5��V�~۔k<R�˝@2��@<�<l��n��NK��ES�:�[�^��	������8:�;����ι�^�tDC}v�;�恈��ح�(��G�I:�g�+���w�9���x;�L����$ !�n1�8Ts�����%*���3���q.�s�v�����N�A��Ԫ5�ԃRɟ�*3%�3�.=����ӻ8�ח{��]P���� �	�����ǹ�B�ȚӤ����t��4�3K��o=0.�D�d����ŷ�ni�Ud7KK��	w>Iw�$`��N���]���s�C%"�T��>1�1�s������K�A4o�m�k��f-�e�R����ШX�F2�H��2��3Ջ�Dp�y�NB�pC�QFMWɝר�|�#��O�E-~���=����^�|��.U�QP�]��&���҇�����=�OH7����  `������2��� F�Zc!��ߎa�Z�NsKJ-CkX������xP憵��VM��{��}��Q�q��R�3PܻYj�|C�9�P�g��ؼ��8��-XTQ^������9�
י�{�NY��p}�lӱ�r��>3�N���@��E���BV)�ퟹh�8�'��&���P0���ݒM�Pl����V��8r��^13�*y�3GCh���D�������KL��A<��
��uү�e�nmE�� �Kӎc���Ő�g��q�2���l��:�@Cma�J�c�fa��:-~h6�N�iF�j�O"u���\��qw��Jx�9�!U�`�j7�<�Q�<�<��YL�-�;��$)L�����\����_�}����\����ܱ�<�(3R���!E�Ӵ1� ]뫣��3!��;�f�ϙ����2�`�~$�'6���u�[9���
iWL�"όa��_�t#�>�,E�8&��&��';� ��P�x�+r7�T/RR��'Y�^D�u�D�@%T8�a�$
��d�U��!���c[[����ꃣ�a}��ZQ�X�T7wC�cK�Y�e�]�a�o.��b#R�G�8�c�r�;��|c��/���a�l#@�J�M�r��J�0+�O�	�q��~�כ��)�*�	����� nɂ��jj�?�*�vu\|brB������a�ǜ�f�B���^R脻�ʣ��|���fO�Q��h>���l��W���0KY��'kL����n*5�NR�a����<_�W��T�ݜ�i���*p~��j�1M�b�,����`���ݤ��o�B��Sv��Z��iqA����Q���c����4���yQ	�i6Kv)�t�����B�`\�$�f>�tW�Ƈ� �W�����!85�VW�CHP��@/j�2<r�#�T��r�_��Ъ�і�F�;vq
�"ࠐ ��~���P����c��F�o�U9���>(������E:MJP��X���|(b��NL��4�TB>؃ۓ7K�P^ukk<F!��}�a�uS8��	�����z��!��tKlrf�W�7ڋ.a��c]��<�]ǜ�M�N}����������]�L
(]��z��4}��^K��	h��-P���L�����Mܛ��@z����N��"Q�[������j��\3��[��T���+� HUg0є�]Z�^��U0?�ל!�4��p�6�l� \���$Zb�uf�8��@e��w�Ftr"�Eg��`�&&��s¼+��x  M�H<�X�K��$u�����5�X&��i0a�f&�4Q�NwB�1���)�� /��,�
�~�٬�m��k��T�!�Z���siܔ9�𧲯>�1�l��8L[,���g�LH��k#�sv���ׂ�;�l��E.	h�4��i�9���3]�+]nmV��a��Ѝ��٘7��I*=3����zMؕ�.�)�F�q����b�./�LFCx5EK����&@cX'M�f���{|����h+0`jn@�ş8��<p��!}�g��n����,�G�b�  ʐ���ƺ��]ߡ�s��EӅ��B_c<��蒠�ۇJG^�"�6$������@�n1���h�k���-�<�����}�����>.�?�
[3�#yj4��W���鞚_�0a��������3�����,u�W�(�@Ӡ����x,�,~l��:8R��z7���4��s�v��{��m|j5L�8�dP=
��]FJ�Ew_��ͤ�����l���ꤧ3�/�4���z��f�B���oȌ���"!��/u|˻B�S��p���M2#��x�δp���n�g���<��ζ�n�1l{T������Q;���ٓ���z��n��r�<	,��G�R��h��r��܁��)��̀)��(��E`�(UK�T��f�Q�wM���Q�,~pw?��6�w<	$-R*�G2�ӳ�m��Nc���<��a�fd#(�Z����'�.ܗ\�9������x2B�T�r���dVN�I�!�qg(``n*�8I����H��AOn�MA|^ژ("��`o�����6��;򢿰w�^h��E�$�	\!du��}�5��b,���� �C���||�R�|ˆ��� c�5g�wl��[e	���.y�4m2�Y�Ì��7"e�ivM�������E��V4Y�k8|���Û��;ʆ*C7�����s��O���*�@F%d͘:���?�-��}F��N%�e���� Z5�����;og�N��'�o��M&c0��� �w�>2�2T9���|Z�X�������|d�q��� ����Kw��j��*�3.:N���x��(mR޼8p��b�M!f+��S\��V�z��~3;�KDt�¤��3��i\�l��u�O�N��[M}�gZ���ʇrS-f�O��*G^;��4g@*#�HPcw��+����c����r�)� ��(�q��*c2{�[�����f�g�5�KI!I�,J}�u�S4����L}C&�zH��T5Y�'�G����Y�Ŕ1��d}�/�����R|��\b�H��ޥ��Of��q��z���9���ú�7��~�c�n£ܫ��[�@)�NǀvD����I�0�
��k��!	�,�w�i�D�0tH���dR�C�zg?��3���{eH�CN�@�4��lu�g�S0@f�B�,4�*�Q(o�u�#bܠ���w�qhp ��dA�{�И�Ң��叇/���U��	O<���y1:��%&Q��\;
�Lr۲�c�n,��"���p��S�H���ձ8���<:��P� V�����^ٯ㻊r7��J��"��(�y����0+��21�Z�^[k�.��?w/�Jnuvܘ}������87��Rz�hiX��6[�_I���p��s�f)IS2#W�o��g�T=����*U1f�'��wYv����n����	zWKлmgc0��YFh�>�_9��  _�5Eo�r���h��J~��f�����4�~*�Ŀb�8 X�/k��e����1_��x���7�?�Mq�;�b�N����["�0]WO����H��`KM\���r���K�bK��J/��������ԉFN&����!Q0���G ��dQ�N�@"x�?��z3�	ϭ��!��b�1`��'ʚ�xňu�������T]`��T���z��ec��p�p�3B�][QL�|���2��ِ�h/�"��P�}�"Lw6�fϑ��Ǎ%�<<L�Y=38�R���R���|��s��8r���{���@�e��x�g�؎/�X�<.��WFL&��F�fوuo')4!e�h� OW��k���ܟ�B �J�lNǉ}�~47@{6Z�tmR�e����D6�����T"S�$x��v�D���B��Y �}Y�E_o�D�G(2���})��f׌�|�I��|1N����ڡ����7�+jVT�[�hR�jY��x}�\�$�0-R������/�E�b_T95!piF\E2�b�Q�0�`���L���%0��KG�f�/`>S����|��$Fc�J+]�C�	��A��g�23�ŋ\L�WM��пN�㲛�-�$�h7�23:Q3���{XN�L'��6{��JN�d$?X3�:j,��0����ZJjιL��R�Zg���p�4�]�i3V���
rr�����U�L�J�G�yE�ql�����o+/�s>�S��6/�T��z�+�h��{]@����[PF�j=��*(=��.im��x��r0�2T������p�ݴ�0Z�����l�p�m��S;v����t�x��{�辵�$�|I2y>d#�<!lO��.����s�o�����$�*t��J2|4I����ϨDҒ��m
�Ҩ���a�^b�>�&���W������<\�Ѡx�E�ޣӌ勺�8���h�^�0{l�/�%�Y�9c++g{�o�l\QܬF&�kĈ�y1ź�A�L� �*��RnU=����� R<�s(߯�mS?�}Z7\���n�5VG|[z0#T0S�U�a?T̟�[Tg7�&��'�Tn5E��eID��{7l���Ʋ�K��K��t ��|�r��K�s��,us�0j�i�1��J���M43$� z�)�<
�B��`̊N6��i��o|3E,#��@|�_�9x(8ͨ��"��7D%�ٚ��6Ժ�6};;q>>mj�"�e�&����H����m��Av.x�Ko�����$P��5cQ��`@o*m�s}�ߕ}���E��u�-%M�Ww��*��e��iv����Y
c�2�n;P�����*�<�a��~�F�:���s���DD%��=D��@J}�e}�y������j,�������Eh$8��"��Ҩ�[���:�HQ!�ఞ�^�a��9��+NN&E��>U.� ]�+�U��i����º�W���
� �J2�UKï ��Eɢ�:.�ҧj_�;7�ƭ� ����k:����T�,@4h��q�j�&*�L�>.���ve��o�j�� �N��~�����Y!�Z�Qu���G�4 +#-����B�5sݠ(�<�͜��dȋ�G�n	�Y���v�*��Y\�ں��.��N"��F�����bƌ���fTwO���j[�liVW��!Xd���y���uY�������K�p�x����\x�Hcg�����#������MI�u�X��ߚW������6=�Y�l�K��h�)��ūfԚex}C� ��T��ǝ!M�ǀ��ڊ�Fa���|����b���Ypl{�k�X���6�x�9(]1�^�o�RrO����(���x7 մr	W��2mP�5k�tB}T�y������ZA-���ui��&g$��O��-����C����-
̜Y��|�/W����[m���C>t.�>E�2:�s�/H1��v�A[V�Y/aG�Ή��(���%|�C�g��;^���Є��6���e�Ȗ�E�\c�7���v�>]��▟�n�+0pqIG&�Fo��4�z�O��TǢ8�N!���yrK!�`�T�J�ފ�*��t�P���6���y/�z^������;�����x�����jS��Y�kW�U�F�Vk���{Q����m��;�U�����1� �/}����������\��9��K�f��s2���-��H	)U�6(͚�x�g0���O��N|k).S��*g������{�dЍYư���%��큄.�# ��%R��egM�<�����ki�s�[�ƌ��_�f�}d�����ƿ� ��}_�Z�燚֌^m>�nvW��%Y��rh�$Si+�(��T�{�)V��x��쟞!uX�-��х�:L�R�[���]�uw�Z?z�L�]_��%����i�l�`����wMq�6?�uGfM���*ʆ�/�ڷ�6n�<4��T��w�����~������ַ��1F�[tL㧥�YY�-�3W�oѝ,[�i��i����3��=�dW�����uE��fӏ���+'~O>L;��;h�1�5G�!�5�i�:Ƌ��cI^:���n�+7i+C���}l�G�/�x�L[�]�M^_U��3,"p�����}rIe'���v�,#����:඙0ֱ�=ͺ��6��t��sܚ��������a��L��O�p>[1�H����L�+��NuG]���u�&�oi�1��t:�=&^𛶂}�F,颼���,3m��m�6j�u�iB��V)a{U�Ռ�AgҠ��8'5A�TF�RA�Y�A嵇��R�8q2*��d�/��1<�n��GL�Q�̌ �D�L��}X5�k�n�u����ӣ��}R~ɹ�<�[�|
yJ�*� %�?�F���~϶��q�������8���+���j�V:IP�/�(k�۱��0�'��Z-_cA��mc9V""�E< m+�c���R�0��d�=
Wa[W鶀���*�*���#t���c[4z�`���o�Mʠ�����f�&�)3tB]�?�+V ˰>��x�⡟F�vR_���)���l,�y=ә���.�4u���n� �L��z�i��ѽ�bjYU�7˶�f��� BӖ���p����r��8甩�B�X�^�����$Q'fE�r!U�����>xЗ��-w��xu�g��}y�p�8oF��<-d��I�rA*���ॾy���|�v8��^[�;JR��ӵ�v�Qo���,��e�V�����nV�����̠!�@WH����R]�
)�A�5�>�q��
�����z?R#K3L�]<�p� �^J8�|��t�,J�f�����t.��]�4�*fx-�+�s������A�ɂM�-綴���'�-�2�GyJ��������kJm.LZ9:�t���x��y���)�Y�%�~K��W�[�� �3�O�;�U�c�EU�[؎�{�j�ݥ̬�
D--�T���*]�\Z����}���z�xz۽��IVh�n�aX<���/?,2�����%yw�D�ǰ�rP��k�M7�o�K��7Aj���V\�̲�����lK
�r��������M��5+�;f�3ݏC͸�;��g{��>��w�y�����腪�U�wf� ӱ��4��0�1?Q1��r-�3���W845�I��K�X��<�-��x�hYu�q/Lܚpy�.�:?��i�-�!^��T�br���g_�b���PI��1w�lPj�D�Д9Q��p���;��������p�a�A�x����co�W�r**�2��1U�	��}�9�ɳc�B�P`=\�<����ٺ�/�y����%Ng����d5�φ�8�H�ތ���7`�U����|�k0���p�k��{���3��x.Q[�sﶩQ���tf�����0Q�|�Y�3]9W�w�q���㿱�o��t�/�>�
~�ka����Zp]'����j�
b��TN_Q��ޅ_��T�F���0ιHk�'M������Aw�2�B�N/s[��{�e8zS�u,N��kFyU0�;-�}�����w�������<V%����k1���U(5O9��dl���P������P%�x�M�U��m(
iɀ7�g�M?�
���i 	�Y�l;�T�~Ec��ȝ�5O�ң��+��>x�_^#�-�2C��B�/_�n���ݾ��LxdV/0]S��˝�*�F�g�t(�Q4X�K�l\-}�͌��9,wi`�Y02K��I$��5��,}>v�m��\J�e�5�E�?"�8P�X�
i/۹�i�4Tl�&�9[�&jc�źn������u�w�����g'��8{�+{jV?�QMMyJZ�~V4۞��63���_Ƙ��d6�X�N`�W��� ��h�:�����nu�V6�O1e���0ÅG-W�I�*-ޞ>SW�Q�f邯��k}-�^N潳\�
)/:�qq�U�I�Թ�)�L���^;���gU��'�&,�j���]=�z˖�5oW�aȝ�QT��̅�Qֶ����3x��ۡ|&�k�gYM���鮐��e��y����*T����>���I��w:AJ'�����M:���aԱ�(Eg�^�7���S�J�u�]6Y�u�2M!����m��/'�(:�t�.���J��?�:h��[O^?��N-7��hS^��|�r�9�_=όg�=�|�������c?,m�_�����f�es^|}�7�>�*���ẟO�\�HܶY}t�����]�A���Cto��_u�7�=,�f�PG_�0�������p[��^ᓎ��YȞtsY��rU���p�Q�'	G����U3?|��rq�j�c�_�����i�W�_|�q��K��{v�I:�?�PP�7�#��ul�,}0e��}���~$sƢ�2֩�5(��a�#�=�|����lO]f-k�{�����\&B��b��SGs!�m�z�����?ͻ�J�.�4���?���j�����a]��X2uS��������!]%�hR��˥���R{�7I��4���l�ג'L�-�q|Z!C(��mWj��ٙlA��X��.j{z�5})�Z3���y�D�F�O]3�'�1't� ئw�������f1(,�⾅�y;5r^�	03�Ƿ��[�Y�KMy�Z~w���0	�;��ke���c�D�X߭��߇�?�B�-H�e��/��NN����#���A׈,Z�U|�l������SZ������Z��`4ï�C3vM��YQ��ٙ����e��9֪_��"9�y��]B�e"��j��J� ��9�`�����o}��P��p�I8��C�Qe ��� ���� ��lvj�p��-��s+����콐�=��ԺfC��~Nl�����Pd1��>��24�QC"��х2yG�~Ua�R�)�s��1��o�O����!Lh�E��B�C��5k%8_���n~[��Дŀ�D#��nJ�'��R<�(����Z��q"M|�>�~ig_a��L�����87D�+R�k{ܶ�o���
C������l�؝*�}�f�lA�.l�U�k�Q�hX�.��k�}ݖVc���W����2�X�����������4[��b*sn����$j�+����*�O�v&�����vya�_�`Q��p�`���Sg[YN�����Ş'����^�;�&[�@�I55��Q�woE#���Z^^����f �}�D9��+�Ȉ�Oxf-��޻v7��7d˵�9p�a�D�����zy=z�W�4D���%QoU�}i/Ϟ�k�#���P��|I�$��	������oJ5�[z�'u|^Z���S��H�T+�Q�����-�َ8Ҋ�RQ���!8�t٥����窊�ʜ#�]�<8��etux%j̓���v
�"�(�����W�v8���[;��Y�-)k��U-���nZ��2�a����ד�vh�؋4ӂ?O��c�-f�����)#���:�<3W���Y�2&c���^RF}?4�X]�y�#�ٵ��ɰ��iw���
�%��� '�-��vҡ�`!�@Qc�����2t�a-¹6��So�4�_\�T+��(��ߝ�^�� �Dz��_�.=�P�a,}Ĝ�F��p�b���Qv	h2:�r�n�[�5��Zߗ#���N:�Z�.uXqE�ߺBC޶G��|u����y��z���ܓ������G�����F5̆��RQSd���Ф�
�(�Z�����$�a�T8�s�I~l�ż^���� x"$����^�6]%Q���o�H��3�Y
��T��2NM��ƶx��,#��Qk��o�]_��G��<�(l ȝϸ 7wA~djH"�b���
�Hxۆ�ݪ��� ��K�G���w��EO�����^�\��6*SGwQ��d-ϑ�Z������]ڒ0ma�������v��H�.Ul���2T��"=���Ŀ�('F�dq������3�A��!٦��#w!�@}�[�M���!.�� eq_U�o��@_t�T�1ר|X��x/p�	�"��<wl	��|����-��`�����n"^p�7��n��{��N3���\x�Ez�yz��ʒހ_���E~�s��I��r`A�&C�{�;�l�f��8��]H^�Ϡ��i^;����M��$��e읮O�'[�����%�/���!�7nbX%Ԍ*+n�����u8@��wu�-�$��	�ɋC��ɈP ��2����Ս�Ӂ|�5Y������7�|�������/C�������r��Zj�-�-rė��"l��hQWQf���Ac���h9I����x�
�vc^��|��Q>Ll��.��Cwjoc!d��<��U5�,j�Do���u�*��w�o�	?`�R�8��*od�
�9�Nh������l��
D<�|:;]�=ͳ;�"	K�<͉ѝ���h�U�@D����\�EE3<���FC,��qS�V��"<U�A���TP�����8��� �k:���=���Nvc���7���\�T`����<z$7G�K:!	3���d]����1o���<{�&�+Y-ԝ~�ٶ���u~n�&�ӦAwսzU�Na���wk��+23���d��V�nq�Gu'��U�rh(��g�h|^�����?	gY�v��smdYK��H9�L��X[���B'z�ޡ:�JXc;����N�c
��T.��nl~u�goz��=gU�Η��̹���7�����!�^S����dKM:���*O�����?�lk�<�1��d�������>�� �цn����Q{i��Y�lM�����]��K�q�6On�s�������B�X�̪͢vtB�>u~N	�S���X�e��p�'�-fz�]�,bء���3`��n�vR���@��Y|�6�P��Ͷ]6���r���n�7����nۙ�H��&젲�3P��R���a�RD���3=,bP��7~��]�C_�?n���'���.���Ho�\uO�\JV�����l�f$�Re��W���ʫ(���O��fN���y}�j>�s5_��`ee&��$88�k��zP��U����i���5���3(N��#-��Ƞ(S��L�|~i
3�>{�,�؄���$:��xQHd���'��>��n�V��l�t�K�$ۻ4����H���޵O�KZ\�� HH ��<��Lدx�&�]2#�-�N�S��8.TS�3U�T�qO�DO8t��P3�.��WI�3���1�f��>I��g�,�"���K�LH"b��������F�9fzY�~����K�^�������ds��⻳�C��u��־��*Y)�Z�5�}�s0s��m���S_�J�����7�-1�@驷�!AV9ɟ5?�ߪ �u|W�_.��5��H�u\
I�33v���q�����Xޟ�ϾL�DY�^��~}�ϧ٩�"��4���m3�8Q�3@GΗq�=�g�gsu�����th�ɣ1x�QVÉ�W��f6����Lk�]gIC�G��\x4>*����y���=f6	��?8��/���w!8|�7��l���p�_q�	G�q��i�\E(�G\�^1I�k��{��v��[���\��僋#R)�����]��Tm����T^�x�`	{��t 2�wg���"�ͷS��#��]J� N5sPT�#g`��H��F��3/���9��O���9[Ɲ��F���Q�;6��,�9�Z��6��*��ww]	1��EG��3C�O���$WL�R,1���y1�v&׍f��y\�;}�i%knj�2noy9t��T7�GY�~jn������G���Ҹ�X�ow(��	�Gc:�I���Uz��p������O�Ti�3b�g���e[��H6R�D^��Ǝh�-M�;)k��f�RE�08��fmZ2��f��ߍ����R��s��f�{<��+.�0�3�xa�լ��B
�����BЙ���&"���J��0'��`�(R06�aH��5�_xK�<7����)�>���JV�3�"3�"���6g����u�nh�Ha�=�R��{t/Ew�����޶�P�b�ꂑ\'����Ӏ�a�d?������!7���g!C��t����I���]�͝c]^}Z�SIM��̈�s2{mwC��wU�Z��0�������N�	w��m]t��u�D��PF�ѱ�	O����d%W��&���N�p����۽^rp��~�
D?�8!��i4�������������; P+/��B-G'ݽ�7�,6���%/>��J�M��e�C�⑸+G1r�0|T�iE��2Y����G�� �)�Ia]��1�p
��fѢ�KS]f���s���7�S��>U�3����b�ܲ|�A�TުJd�΄ :�����Z����6���~��54F���}U���9�엉T���Ǝ�w�pYՖ����sx��j#�ϯ$:L�u���`�vr�tx'A���ʣ"]��t%�����=�z��aۭ��ڌ@E��_O�(4r�*Spܩ*&]+���)s^�cXQϐ�id�2����(U0�B�va��=�i�1y��\Z�&c�Li��*d"'@�<�`\�>�_|���� ���R���q���z�q�{R���6��еy\�Q�1�̑%��K+�N�ܼ��L_�?�=��}-zi,=�b��.[���b?'II:OI;��3߄�Kd�H �B���-g�xP�vD-[�羁����.Z���7��:�٥
b8q���3x��V��`��K����r�|�V�9��R�q ��WE�ґF0θs}��+^{a�F���%�o2}��ȣ`�5��5z+@D��0�N�~pK��Ao`T�R�AM ��k*��oF{�����,�T���m6Z�<�*��`gά5n��|&^60�3ʻ-I�2�7%��&�x�/�}�6��!D���K6��$B�g�9!l�U���Ed6e���87j�錈�i�^\�ڝJ&�I����O(�tc$gߵN���ئ�l�pu�.�*bH,�`�D��B�P�N:��Z2p�G̊:���r��on�*D����3݂v��擨�C,�DM3U��Ls���9�2�Q[9���/q_Zap3{Z��j��.����w����ɜ#���Wȫs�gHn�/�����iz����������Fq�E�s�.TQ%Cփ��D����!Ag��v5����Ą�hS��1��V�D��\ev[lU�ǈ.*h�+k�R[�Bw��,��:�ie(}���>"k���W���mq��~��6*C�^���W���v��I�|�R��;k�|��y��������MX��m�:�3�#JetiJ��O��G��z�C��s7�>��!��t��iW/�8��@����G즴a�����Qz����*�x�[�kx~USٟ!���2n�֖*4"��_����A��]Q1h��\�MV-4jJn��jR.+3ݵu}��KN��y[~U�vŸ��v�6Qv���]Ň��_Nb]y��!~)�<��y/7���VAqT��}VU>�����/����Mk��o�`��F�?� ��j���b_�)}�����#��d�-�����*����#W��D^���s[���~�����N\�3����G�����f����o}w�#�y�h����{�e�{�6�1�TS-:�e:|p�{�Xho���r2�4W����`}�OR<���`D��؋�}v�߳�?�L��٫����[pM��17����&������&���d�bN,�����_dK�C��`�0>ů��֨� R;K��ͧ�w����4l�,��t%e�ӽy)\������}s<�bp��~Y��?��y�9�����1FI'>���o��ϴ�  X��B�oVI���+l�ҷ���;z��!?�vL��G��'��F���tSL���9�����߁��^�L8�u�;y���R�?9�dR��t�B�sn>��7k�}{�{�pW���������1���Q����IH���P?��G%g*��r�d����ʽnu�gk���z��Yp�lƨ_��7릭��۝�Ĭ�%g����(��e��5m)"�d�WJ!�+E�s(�·xR�_S�5���wQ���Q�bJa�B���И�u<�[
"�n��9��\��[�7��>#15e�hm�b��v���(n�Q����x��4��e��<D�EUEቩx[5F9�e���ā���Au\`EQ��+.����_����)�����\�1'1S��Xwz6��3���-f'�?=�F�>�%�����n~�8���y��*>%G�V8\�*f�s�����1��qk�k;�n��6�G��k����6��w��:S'�4���lFw�	���۱W��Y9.�� ~��oIœw�	yF|t;;K�;���)t�jM�:hAp���G�=�P`�-(���/��E�{�}�*z��Ҟ�P�:��B�pr��&�����ɣ�'�n"�d���iB���טE�5����N�؁��-Y�����;�a��n�o�*N[��љX��>�y�MX7�$��w v��
�	������Z
ɜa??���<���ʦi�y�bAaHu��Rj�YI��J�EC�ǀ���ܼU��>4&;8����ޖ�w9_�L�!�&8H�����1�$b���h�G�.�?��&��\l�zq�����T���iH������o�#U�2I�b�ѥ�.�b��\I\����������J}y�0��s6x��}r<�=BL�r���]Y!����=�\'<?@xޞ�ǧ�ȗ�Mfε\��9�'��KJ�u'��C%@W�!���:qJ@�Tz�wN.�L޿� Y���V�
\��{Ԗ��Qr�K�=3o���f�ef�=`��>�l9�
a��C�E˂��-p���G"���Q*i�[νc����[~�E���W��5v����&�k����k�b4�)�ʣ��w'��X�������e�9�R�<=[�����	��ݾQ
��>w��ԣJ���e��;rtB����pq�����x�Ym�me�b 9;�n�	�滿 ��Kr�h�����`#�|C*�Q�]���+@����Kt���DUGU{
���[u�^�ܣt.��F�Q&�,��LUy�
5�Q�6��!�z�A�BK�=���IۆL��N�8� g�_�w?/q|��[�kgZd���o����(��_Juר4<��W/�0�-�3� 'rڝN��ˮv��,R�ׇ��C|B�x}⏞_�'G����>�r��?	���L��t$�X�wv��>��Rbq�����"��4�3�T��R�u��ӱM�|�=�l��$�
^p��H���z˿���x�B�e���{�B���o�d�Vh�)k��X*
�fؾ��.�D_�7J�O���**t�E�K�?]���avT����0���l{W���7u�B�����F}x9��c}�:w�����U��&(�TW;t ����N`�Z�gC7��ʣ�9����y{r�z���4�)���ʸ�;�Ya�Ϲ�ޗ
�;+�Í��lG�?��7��嬫(��6�4���	az��o�pXKH��iu�ד��פ��e1�潤�������5�d}"E"�z6D�7�����x������t��D��^2��y�^Nc���X](P���qd����"O��Z=O�_�OU@+rp]�㌷�X@Su�o2�����u�r�A��@0H�� Ɔ5}�[�2�Tn�dnl}2Y��9�뗱����.�WOĹ�e���㑻Ri��]�&��%��o%�Vau�-|�_�?<�kN�]=�'�B��q�2��Z&g{��se���ȂcɈ#l�Y�a�څ>�+��v��ma����3\�m�\�����D9����s0������HMj�u���XD���r��t��,�����|�,�����:�����1ݴ��7_����E�&#��^�bB�~q��n����(t�\S�Q�W�UO[��pw+��!lԗ��ܶ�5`A����Se�k��)O��l�V�`��x�ɭmĨ`�셭MOI�Rg^.��!��4�A�w���]eUJ}���.�x���k)��Q��GA|a~����R����޻��)�F�5a���U:�^EK�^�3���-JJ,��[�t��;U��I~o	7�X �[c���ѻ�WQ�6۬:��S]\�J��e�}�zLG����(�ܥ��*}b�)��h+_hd>
@��H��f	&�̹�c��!�G�(v�I/��|�Qa���n��V7m���dEx�^R୸��h��Z�\���R�9$/}�4��.j��hd�ҭ��bj��*��N���)`_'��3��hԢ=��.�
��c��M�X���Y�M1,��Ջ�>t_f���/�v���K��[�"W/p���V�8�B��wӮw���
+Q�;�\i�1�;k�������K� 4�波���]����(��c�����>N[��Np�=�ˈבt�xF>T<ƅ�O�`��ð��R����\�F��ga���('`qb��a����*�z�Y�*Q����Q��2&������꫒��V��xu0�ݫny�)�r��h������FH���]���]�4�[� �	�gۜ�T�[�Ky8M��v��߂]�>��0��[�HU�m�Մ�e7�B���#��ּ��E���^tBd��e�󭄈��P`G����I������b�BQ�g�|[ܰ�Ǚ)�X.	>�W�6b�����ڮ����q��[9���S|��@��Uř� �U�H�yD"s�ii��R�݇wA�G!�o\h�7�=�G)�}�;y�L��8��YVh,�%Jw�{��EƄ����X���.>�E@���fh8�U�S#/���בI�c����MDN��/�%��Y���[t~��%�h9yw>&Ŷ�Fd_��)T
�M+�V\�&�@7i@�L1O����5O�Ό�����:���[j�ǍÛE�Owdަ�5,ݤC��tL����)c��FģA�<GuRU�J���� 2��Qګ1�d/�����*�sRֲb�Vw���Q��(�/𽍣V�{�9Ȣ����d@w�ہ����1O��1XP8j���Wu�Œ���QNdBC��������u�f��]mF�Yyc���`.�S���4AӖWv6�m�;�n��߰1�ǫ5�ɗ�13m~*] #>:���hmY����R��4�Ϲ�{(���
��X�/����s9[lŌ��?��8�Gܓ�,��{�����kݫ�E[�һ�
�_Y��w\]$�)�VbG��\�b�M���nyl~#/��u%�(Q�#�Bjx�&��vQf�b�/���y�)�p�aP3�C�0�")�����;��eB�Qz�;Ύ��^�k �s��+�s��?԰�\���{m��
���v|7U�r��9���F1I���볳~K$����Ѽ�d:�	y��5�]K��R�	Ai8�������t�L)t>���N`$�#�KS/[1��0Z���i!%ݴ�r���p+.!�.�hG�o�mʷH�0���H?�R0���i����>}��Q+��-H�6�1���9P"������_̾F5�@T�N����ˆ�n��5�~�8�ux{�ܘ�������۶�b��H0j�u�x�|��e�������G��S.1)ި��I�ū8�z�P��\��o���&��T8���fY��M��f��=�U�Ex�A�]_�Q�����Kbp8�g�bM\'A+p,���q���8�F�A�W����7�DR'��줝��r:�E:�C5���ٮ��xJ��= $
_)���>
Z��Ѷe�/XT�a�u^�b;e�wdO{^}f���!�aM5�L����+�:g{����~�C��׬�/�}�M�+oMʚV&�h$��. dM"�BPa��~��'������m3���3�5K�(��'���d��6�����ebr^����xr$��[r8�_���3,�8�xĤ������-��O\����1Br���>�s�L`���A}��yS����"E��ILKI]l�6�E��h'r��~�2ttQ�����
E�Y�x�qmY��?�a���%9x��cO��(��(\�=w��Y���t���8���N
, �f
0+��s��itZ��}��m]{ľ;�z��z�w�@|ǅ�z����_�|8}ZgOo�;ж���.uJ-�9Mh�H�މf�Ӈ�FVR��ǩ��t�~X _ߐ���� ����M��n�÷ط�ang$��5��]�˫���W�tޱͩlRw�T�GG�di`[l��l۱�r��c�:5P[n1�K�G�,�0_�-0��F�z��	�T4�s����[̲���{�S%����+�;¢��&u�]��I"S�PZ�г9��N�]=z�]��؂u�p+s<�vRЅ����2��w���1�?J���*�������{��m�;+Xdk�}"L�&�Z��s��G���#�
Y��B����J�*;��lǆ#a�0}t���+�d�U�3A��g��V����xg�'m��b|�A�k�n���2�� ���/���ԥl�η�DYF�ۣG�(��4�FY0�($v�s�A:�g��;Ŏ����[������
��>'��@��+�/`tT����CR���&D[-,�\)�|u�\����e7lq�K��Y�V{/��=��8|�3��������.����P��^rvOߏh��Ca(�_ɪ�M�p��O�P�/���O�@�{j�z�a�pb���zP���\�"�#|�B�6��N�-�
%�)��|�֪��R���3��Y�����5�rR{�o���'�9<����W}� ��$�)��#��#��SO�k�V/�GcM�t�=�4�v�ށ@�L�G�%�K��x�E��"S�E�zܙ���q_�_�����g
Vw�M�(O�fT��p:����qJ�>�q�;���9deP��W~ %!9��������%���m��?\.)�5�/��hTS+?�ʓ������R5/s���;�T��t�7xf����lT���h�]+�c�r����ѬBk��5=,m�p�c]A
�ө��_Q�FNwn��k�%8�<������҄���Q�����z[R��ǋ�ӎ?CDJ�/��À=;��o���DJ���?�0CCq��0}n��$8���G���s�8�x��c��M�,�mӎ���:tt�;������4���N��.��#��:*ӊ?�=�LS+�wfE�13�0m����^B�����$�z�$�6v�F�-�D��z����7��C�H R��l���R6i�;���鬜����O�w��[��}�	wd��k�֦��ԓ��^��^?Վ�8z�#Y-�v4�*�w)��2}^n�A؉񧯟�¸_�~�ö�d\�>_�sɌ�ɫ�_lr^����޹�Sug�����	����RX�O-�(U9[I�|׼v����J�ì�j���炞���!�D=�ƕ��+�j2 S
�VH^}#gZ>��S%�9܎�W���>��6[��@O*�����춊��`�T����Ě�r���[���5�e�]Eف, v	�����t#�[#�fVM������6�1�	\pS-�	C56�V�#^u��{\v.p��Q`$�1<�sh�A�0�@d��:+E*��eƈ`Z��^��$�&��M�'k�{{$�>������,p�%�h�qڊ���<;ۊc|���8�N��2�FF!�xH��l>�L�Q9$9@�ٸ��S��{;��I��?�a�s��np-''}�;�Y<�~~t������ T`�|T���td4uy[pm*��Zr9g�g�d��O&;����/.���g{
����p����^��+��/v�DɤZ~���G�[]_����z@�i�wRF6L�)�ܫ-u��Ҳ��-?�w��ξe��z�Պ(�8�3q�bs��m���cd4!b�axvdW������6���L�!mm���Z��`���o̶Bxs�;�8��J��w23q��t^$֫��G�y��U,p�1e��"�X��(Zx�j���E�(�CnD���N��ę���-�	YvGUZ�HR�Q��Q<�}�M袀�3vWJ�S��T�ң�1���c��o��h�$"�]�N�sH��!Rx�Ng����=�L�N���"8��I�w�C�Ww ���D��|X �}�(�їP��ܓ�X�8V'Q&B��d���M��Y��4u	�K묽1�)��L��U���R0��V����)Q& :���1�cφsB�`�D�j�F�nQ�^�ۭ�c`p���x�l2���:���
�Bx Fd��z������s�T��๱�O��>�Y	����dq)�lI������H8�L��Bg�n��ؾGף�HaB��x1R��B],��=;*6C�ZL�R���'�8r�)���d��0K���{�Jn��5<27�!Կ���>�}%ꠀ��
T�o���o�k�Y���|�C�fҖs��U���O�fG0H�E��lG�8ݦ+�3�7l-�`Ҟ�Xb������\A�����������iǄ|����¥h��ImUՋ4x��W�\�~Be�#+�Mڛ39��:�~�,�H�����y�w�k�W�����,��YӆicS�ᤣU<L�u�yUA��?"纠���7�ة��iR�h�����.�4����Ch4��ҡW�7s��"��T;�Úx"��J���l�F'<�1}ُ/(@�=���6�T�j�����6C��%�D<��e47_�X�������19Ӄ����Н��V�A�$f�u2*�T�8������XT,���m��|�/�M�0!͉N<�@���2t)�5[�!u�e����bp�X���{ƪ���ƾT���{0K;�;"%=C��J��J�zj;s2Lj��c�A��6$H-�+U��6^�"Z!1إ�-���i$�����+,��[#	�;|�x0蜓��{��.���|��]�ivI�^���������P��`��Jz��ll�]�HJޗ���$]�Ǟ�*�W��Ʋ��} ��Ș���z᜔*=�a��m����ά�����J��0��}_�5RX���/��U��O\��⽊�c���&d~B��B�p���v�-���p��e�q��:�Lt�.�m�����D�]�sv���7��[��!S�Q�a
�N9q�v��!;�ʎ�uI٬V]cXr�3����Rw���f;b�.�׿>E�����N�F�C Λ*��11p ��ș$~l�V�v�-���H�
����Sl���юg_>)�~��`a|~qJI.K�K!=������;"?���xV^kT��؈�ݜY�5�;[�8�a]:�㢶��� _�����JS��gb�eH�o��=�5�g<w| ���cםyMg� bE�;S�}2��\j-Z��"������U��?7u������+J����o**�-w~�f;�l��	���[=��I}�����X���3���~i��E$��X~���7��!�# ��j){�u���sX���%�!\ӧ2�|�F~�3�n�4��v	�("on��&�p�y�&�3�Ű
G����@[�7e��v����/����y8�\.�̥���Z\�ZX�ZD��8�Ck7I�Tc�MU��HN��GP&8���t�=���'�*x.]�4�:
.�2h��G�\V�P�T&�n��F���wb��><�zK$[wn������9N#R4�S�og���R�1�S�����} {�)��BT{iF�F����?��'4�Y1]T���*7O>l�QX��ػ�S
�03^PwB�������k�V��I�� ����X}�.�t�$*^�}�'Gv~�䄤���5�RE�R:���������1�
DO,5�����8���#��B�<�lP[L��5O�o�Q�C� �ƭ���kiCMg������L��vV��=�a�Dt�$m��w���'k�6ϸ����֔�Xa���K5uOB���ϚH)i^L{Z ��qiZ�C{'��}-�L�� =�w��?s���v�K'b��pq�V�z<�K�OX�7�@�.�ݾ����|��g�,nl�nz��O�x�T��z����R��P�P�20M���"(��KZ��A|I����F�Uhg��c�=��S.R>ߑK�W�
-���jB���tV�F��]�����06�rs�,�4�� ���Q*�"�ð�����&۷}ii	IEJAB��!  �"--c��)�)���T�F��F��������������<��8�nV�:^0�ɵ�Ts~& I�K�R�]�أ��x ��А�:� o�~��uQ�{y�Q�tda�H�l�ɺɐ4l`���,"��FQ�%M��O��Z����, Q,�M���;�1�} 9�vlXA>
�1����9w�gD1'P��w|tk�I��F��+-\�˽����������.�Mg"�c	,*wW�3�h6qF�Ye���+�(��G�k#?�)l��
y �	ٙ,�<UOX������k~pB�f]& &sM}�	rZM[�ge���F���	�U�$	,�c*���"�u�~D�e��%}�P���N�k���ɬO4���s6�����TçC��%
������zCk&���Qյ����y��B��l P���_��5�a�7��+|�IE�`�ÇS3,h(�JP��u���B�_��^9.]�?4딊nߒyד�&ڸ4���NGN6���l0�=K��.Vr�u��_ֺr��C,�f�;���'Z�2�RbIP��},�ꑤ^��X���S�Nx=t�����C�/�*(�K���t�dX�5w�m�qQw�Z� �n�̭ͫ�"�qH�|��l-x�q�;Y}�|�}ث�&����<�_� �	r�Z9�����,|JY����^���G��\c:��?+-�����9<j|xז�N���`_��5�4Fpу�ۃe�y��l����ߨ�F�;�tfD��|�Jri������w_��>�A�]�V�љ1��H0'|��4���b/�ok�ؔ�Rֺ�?���K2jx�e��У�՚�4ҫg����g@���l�O�^4�텩\3�7�����N�'�9�����O��`�ZqT�[@�K1?�t�8�&��=���<���G���8�
,��T��c��`Sԥq����:�<�޽���#C��]h���em����a���q���@q�J��%�e��D�6-�UkkW��`ZU��?G"b^��*��ڤ�Ds:���L���w�&{�v�j��@<��T��,N����R>|�\�����$+�#�c���0��ǧ����7���q�In��{�k �?reT�®wƲ��zx�Ԏ5�Z�O�\y��:����g�[V,{�(N_)v�@���ya��VŌ4��DS.�;I�	 ���	i�������S)�YJ9^-��X�T���=�*�����J��q�YYK0;}��+Q7:�2b`]�В?C����0�|��)�|�}���Ns��]��YR��R�w7e�}��Ѻ
��0<X�f6��tͯ(Y�>ʴ+�������x�e�;$C"��Z�#�]L?_��hu�f��!c��Oi�Ӓ����W*�����n��w�R�ߒ�[W�G�6ܐ�|�\:������?�cs��i%y��z�����W�o�j�&����O$k([Z�O��w���������`f���rg��Y ��Q���QT���F�y��f�Sn6�(Il�`����Je��8�
�ݛe_�[��R���CG�F}S�3@��GF!�#��L\=��������z�l�fyr~鲱��o�Ӭ+y�@d<�}�gm�H\OC6Fe[�x�@�ʭ|�$�浝���l�lW�������";ֳ��)���[��p�}���"o���ҭg�bM9Ae>څ���gz=���t:Χ;�� 3�Lm��\��1�>�Fl;k����ېS��?�Ҕ��L�P�l�IF� (���|[=���-�D�I��E�_Y%���sG3���4&Tc	\�Bg�$�ӺÐ(3�'�e5�����g78e��_pQ\�E9�[��Z��>{ujq��O?�;Q+���xPO����[�@�R�0[`s��%�ʳ�gԚ#��L�?�3)�NL,��d�!3iY1�8e� ���X�>��Yw�,��?�~g"����\�ˣU,��7��@�9��+<y�FO��]�b���P�����bj_��7�
�Egׯ!�8.ܾ�bŤ�7^-�,�/~ufkt��Ʌɴd��mX�=���&�nvL�]?�A:%�ƥ��,Q�ϥm,�c惖k�B���|TW$9�����_���NiF~���O���i*^��5�����/����C�D�$�wk[����6n����D�ϴ�r�� 8李�o��u�
��i9"�G�7;���o!}�-�?�G?�\��g�X�Q�u�3�DԂ�W[���}X�k�tv���h������rJ�����]��L�ڧ�M��:�ҰW#��ɀ���x;+�,�X�#�_��_?&��1�  ^Yo��
�_Y[����=�����lX�#Re��@m+�ގ�/�y����E�x$W���7<�RU��%�&���y �j�2����� �,�>���M�r��8���2yB&��,6���|�R?���x}�L��T�3c���I�2�ye1Ҭ��ї�M��s�4�ּ�a�]����/ѣ���訨T��6���c"oa��C��f�,��h��� pp�$��8�;w
�*OX/��\vkko��'ߎ*�]dZ$=�&�����yޞM��GX�䤒`�5��\;Hޕh������*�Y�?��^	�	3�MOz=�=���*�l�4/�E �AaX��-d\�k:QBF�͛�?i���/��s��_�Ar�N� M .jzU�8��ʏnԤ�"�G$�9|��|l��:>r����%-�k���Y ���`t��KMm���~�=84��Y��O������P{�b��"3����O22�ml�;4y�ꊦ�;bے��ߍ<X����^�s��f�Z~�1�����c��A���6��5et�w[~�����~���׳<Fۆj�]�:��N^���;��߄ضS�;:�Ʌ�	]r	���Nt;pRc�Z��oIɇ�X\��~p�z٠l��,�ip��<�Zz�����KP߭*�uȕ�������z��'}�JU����>��.� �U�Iy�k>]@�IS��~]s�(���g?L^�J���<�0S4iͻ��Fێb�
�ޭl?c�38;u/
�(J�1���n��O+�����G�B)5C})u�qj`�L*�P�rF��{��x�Wr��*�9?����}�;vӅ��$$���(,E�w������~ا�$w����?'])Z�U�Y��LkW=2����ޮ;�e+jV���q���/PY����S�l5���6Z#T�q�J^Z���4^�]^~j����B"3������O�4�ͰKm����1�~��P��ó�x{�����z��Y?N���`���P��ݿ[����ߊ�ډ;��]��%��}
��~?X;��a�;�uT��塀����}����ebp��N���G2��I7=�^�!W��gB��+VňV�ɯ�1�|���?�	̕R:	���X?�[�t�nl�eiN��	dd�ۃY���*����q`��E�3��Uf�� B�.ߺB��_=��;��Ԇ/_
�j32ķ3̛�f8�v/:�Q�t�}vBUe�2���v����V�&����9�����. ]O�k���mw*�Η���IU�&0����C�����OM�y�g͛���WY[��(~����']E�>qa��'��2m��F�SS�/Ь����Ш2�*}n��z��[��Ip�Z��"�c��@�,}O� b�0ِ��C��ã�F�� F/z�X�rL(�4��١G�����̒���/"��q0����zب�6�&�hB�_f`��ӧ	��e��#ѥF�9���� M{K����h���ζ���<�4v���J�5�|��*���6��}����+�5����|�mf���z�r���������[ڟTcLR���ƚ ?�af�m�қȤ}7/�o��	�����/���]\p4��o$��������$���}��Y���Ύ��1�F�4���Vl&&�ap�*����S�Y^�@�U/(v�%�)��A����ی��U���<Wx?��1C"a|��<�n�r�� �X�F�[�b�u�V��_��-���Fų�9`֚�,�îj,��j��x6<�|s���{�M ��⤿匞����}�6c*��`1L�nv�"�Um�.�L<� ��hM]�m}4�����eh�4�/݅�gm��˛0=)/š�͈vG{6�a��ie]A�L��iT&��wf�zdM�[v��|7)A�A�W�GV
��m�
�kvm��y��[�\W�5=�%�"��xrDy� D=�9�ב�i��ݸ>�dJ6�:H�7V*Mաhq�����v��n�z1�7�^	q1 �k�_�ҕ��I27�*9כ��:��qְi�`,�箄6�Cz�K�#>��C��(r�*��W������Q�E*ܑ{w����5�m#��l��"�C {�L$¢�Jf�+Q�?�ܑ\$����W<h������[�����a��!�������(/�&���_k�k���i�v��`�J�T��H^�t�<�+��a�H L�	�A��J-��ӄwar����(�q���]��&E��U����D|���89)�I�2�~�v�y��\<��_��5��n�[��9bB���彿`�Mn��ׯl����� ����lp�߶ɷz���|���7R=�B'y����fq��^�1t�
�)j�V��I(d�9���$5��ː�+��
��i��6"�����T����u����\�>��l��Ȃb��#�%���$�WW޺���\M]򰻷�͉J#�J�d�����\�����E�Q��v��.�W����y�7����2o8���p�x������:D�_� ��!�����w�n"����M�껓n*�k�|��kð,ЬQJ7���|�����O;�B��z�7�r���,Sr=���Ն�4�ՕOϝу{35 �#��6�뤔�Xw��/Z=�Cu-��7���������"��?��������B�Td��v������۴�׫V�S`!�` _�v~�U�\��pyYpF���(l�����`�>:���߳��k�����^s;`�:�>e�Gɛ����/my����_��|f�3,����k,�y>�n9>����U�]݈�X�f�X�1��T%�HX,��>�+g��$����>�6^�#n���"�c�����m�j��cmB�b��E;�t�}���©�_�E�y���Ml;�^���o�3p��+�xµ����ћ���'Y/Y����+\�+���F�8��Z�ޡ�H��B����Qw� ��	55u7��jѮ���4���������D_z�c�-ġ9JW�K��|Hdg����{2F0&�)�\��'&�&C��M���;c��Hg(FE�3��#p�<�嗯���b��6�)R9�/�`4\Ս��a��ğ���Y�ǎ�?R\��&2h~ﶔ$㵛D������p�*m�P��_���"_�Q@]O/��ծ�$�Y�%����yN�0\~~RR~�i8q��{��i�:�F׏P	\K�Ϻ���M=Nnҝ:��ޑqf?������D�{����&���R� o-�ln��+�ƧT�^rՃ�cZ��f���-甛'�d)����͙����3��K���u��?��3D��Ͼ�����+�#YӉ��A7�v����Z3����9�a�&���]�oI�_���� PA��0(X,eD�����+i���� y���I�f�1��5��2������ ��@�oG���#�W���D�o6��0�ν|�;�������a���1��ٚa����k���w�3���~V�d=� NIn�uS�y��>��\�;����o$�IxJ�."�ODgH2�@1d�-+e��Y1���8�h+�\��=�:y��޷���G��V֖�Gǋ�qQ��i�+�(��N��R���1_�����(+��ֺeK�'�pUmmNm����t���%�W��U����tn��Ug� �gdy_��Ӟ����q��e���!fq�G~7��T����x]���/W5�8��l���"r����L97�l6�L��	ʭj�&�Z�{�u	��.)�!P��݁�l�6�A���+L��ٟ[%V��\ؐ�L�ϵւ֬��n�,��<T�}2� ^�^|�!��]LQfQ��}ݽjzm=�U�@B��F���v\����dO�bB�	�ё�{k#��!�<���64�}^v�ǜ�[��{zJ�2��Q�􇏓�Gh�������7�q_ ��#Yv�w�R7֝?���/��|_>n60o�����:'m������5|��0��:L����q7;s�?{�v��:R��y��#���i]�U�"���!5�����q��V�沦��j���kq2PM5���+��{=u��3���h�)��Ȯ��
B�[��Y�}I���@_�������̟�A9�/߱L���'\���m�ζ1��)�͸^�m���?�H	�l�ƿ��S!��(ptW �e�|����|AA�2�H�w�R��.)�V��S��ɥ���"�_ߋ���_`�H�V�-��w�ԩ�Q,WY����1"-A�,_�qoT+8e>�Qw*N=�a�ʬ�ҋ���"��Ou���"�J�F��Qc��xsz�_����
�E!Ќc���ɢl������y꾈�Jt���ES5�o*~�Ω�mq��C�}~5{��y�ڹc�ݘ��(N�x��mF�ۥc~�Dt����8�����9�A�1�k8�M�y����cd�UǍuP`s����vO4�h{�X�!ׇ�'�=W��]T�T�b�_�l��hɀIE�O��0	d���)�	�'rO�����>p#F���ӫ��\��ʌ���z� Zt��Κ| �dR�����=q�� TU�Y��jk7��F��w���%�U�T�\T�ՠ��pץ�"�H
�Qb�73�W0Aa��ɑ�g;�E�?�94w�r���.![7���81ݜ��y�;D^��@1D�qSD��;y�P���A b�e��z^ѹ�9�AJ��4��jm��Ӽ��s�}�X�/��6w�1u6��3�-��������:�hj[��8#ӥ2r��E�G�;_�:n�v5�Y�ב"xI�"Qڊ
���� �=Wܬ��|�פ���G��:�C�W�|�/B�d�
��l���n��E�S_dL�E-�L~�h���,�����A�p`kzM	�=�q��89�m͡��݊��1��j��2�����,�����7��E r�տ�������s&Q�;�O�0]�n�c����q�LL�,�NUV���{إ����V�_��ZE�a>�8�5��8ͯ9�D�G��2l!(-�Ё�T{j�V@h��Zdd�	"��+�z����h���ac��;��Q�O�Mza:b�u�@�:N/�c�ne��,#ƖB���C��H c��S��H!�8R��o�	h�Ao�5��J�z3��~G��~�*U�3����nv(k^ow�̄��/���_��ˏ���q���ǵb�ٻ<��A���F�6Zc}+ߔ�f�z��`D�E�39�hԓ`��ܹ�N�t�u�7��d~&��R�}*տ9J����-_���6���5�l�;7��XI�t���.�^��ѡ�JXj�/����m��@}�1�<d�X{"%8���rz���)"�ʙMt͞F���H듉��t"�1�{0��w����s{
�T�E�"f±S��DNt�V�M�X}L���Ͻ��.���<0T�����l��~ILH���� �TdEq߾����Ddo��ޫoceGb.�`�`0Hp�0��*D��"r�fZ2+�h�u�ୟ�}B�"��CN���ˀ#!J9����^���W��O�61�"{DX�	t����+yɀ�h��V���h�{Z����AM{ϫ/��=@�ay��0=(M-i�<���k�zR��_�%��U�F��w���]�{K3xE��*z��˰rØ���UT#��!�7�/���ڜ�s=i��%�K( Ȩ�=eQ�؏���/E�ҳ���7����J�8�C��<��w@�C���ߴ{=����g�	���g�2<�����j���~Nr�Q��2�zů��`.���]�Q�l�ц���X��	�G�>���دz��O��b�n���ר+Wna�]���rv��'m+K*2­�JxU�'ș�,A�)�Ҙ���8L���FI�ʚ&2q���k��e�X�due��	ud��G�P�\llx�{�Ō����$�z㣫a�֊��s��ɽ�z>��!�����;-��v~ƌ�5n>�A��#+�ס��c��<���y�Ql�%4O0R)L#���1m����p��[ېڸ��SGZ�̼�;��QJiq0�{�{t��m��ki���z	�_>_�k@�X*R>?p�;��}�� F����aVXP �H��z$a �B�ňyi)j�z|��ϩg��ؖ����p륝3�dߥO�8�܆���>L*�z*VUX�SR�%���d��쬣x�u�VY�	ɣ����A��^$��c5'���U�ܒ�6N����z��G�m�u,�碵:��V����2�4%�#Պ?�d�"�L0h5ߜf�%kd@��^<������奸�Ờ-����T�����ۈ��XZOw
{:#1x��^	_�$��FK�6��=CZP:�7L��>�g�
o��'�׿���1����ɫ��2ƙ`:�=��H�<�XG���>P��h�<��hU�8^��P���3r����2��{��T��;SElm�l(��#� �@g���לn~�c������櫡��V�r!G��Ce����]����%u�0��x��&��s���w�e�lOUj�yø���FQW�ǷDS��_���r�;�5��QU&_�6�p�IU����Y���T���2���:��mgw�a�JL�=a���c�����ѷ&��T��������>����ؙ��'�#􂫼z��C6���j�:�u�$��:��t{�j(Y��c�wJl�ךB:β;0:tX�Z;Î�f�9�Cy,-��3�����*�y�Y���Ɉ|���|UQ��f��\z�z��&�����jģ
ʛ��ȩ��7ϴ
�QZi��k���),��(�
#�mJ_mx�7�ƫ���S�����)i'ڤ6��#X��,mx�w7~�1���l�5x���漗��=��Z/@����}T?d�;����J�-����^�'�?�?<�R�f8�ǾC�-=���D�e�8�����X�)ș�2SЈ��I\}F,lU���~P���	6v���G9Yk@��?/�+�]����8qR��?Kx����8�{Q��߂.��^�PQQ�s��Cbޕj���G�t�	:��zK�,G�P%����� �Y��]����!�?�ȁ'����a�MpHe��H��k�Nd���@�+���G���7������!-M�_����s��1����b�4��(�!�Z�_n��X'� ���~���һ�f:ǖ������i��Os����!���#�>T���k�0�P��Ra()y	1��'i��a��t�n=�[����������gͥ�oݟ��B�0����A�[�0NL��U4zx�@%�l�E�WT�W����v��S�L1;@��$x���i]��}c�N@�="�b����{E��蕃����=m=
���K}��X�g�Җ�6�;ƞ~��^��+(d�O�����닳}���6OP-�2b�2�ҵ+z�Ȁ�:�l��`+K�"��߉��l��b�	�c���-�uF��'M����X����L��s�o��й�
�.�_��C�=��מ]��g�#�#���\���ي%����K4�*>�e*m3_���9�ޅL6�E	�ba�K[[���:����􃢨��������߽ɸ(���\����ޗ�&��:q�z�D=@����%�QD�T�yk`<�f8:0�
~�(���������>0r�tG��rX8�h$y��I�Ou�S�� �8�������*�U�@�5�_�X�$N���[��Fļ;�z"x���G�#�p
MK�̰���Yb0��;|�F��dMĂ�F��K�ڟ�O�fE��i=&ٴ�������s����ʩ�e^չ�]q
o���u�f����]�bu���f_��S'.X�t����9����**P+�F9&p|?�RQj<���S���(� ٸ��ϟ9�9y��C��4w��XY��F�ߕ��� ��X)��4���Ы>^>�"���TF��#<����.ٛ.�:L�fRo��c��8��'ġtB:��<�Y�oWL�{�t.��p�=#��L�@~ �t�c����3X+ړ����Q�l���8��L��}�@��_&秒o�TP��X ���m���L��NGmJqm4R�5K� �S��N�3DJ���n�P�h�6�5�m�p�Z���cꔥ�c�����y~��q�v����>J��9�@���kM�����k�݅�X:�?e6��a���o囱x~��#��RE�F&�<r��k���H�ls��.����!k%�h�='`�B����;�h+���s�l�Z�Ş�Ĺ�+��jȟ�9���`��Ł^Ƙ�۫pQ�#�%u)�>q�%��9��D�9�f8'���M�MD�<�:ۭ����$�.-�u�Ap�ݤ+[�`J⛧��*��}F��eD�ëf�uo ^��9`���öa��gt�a�]w�n�;>����N�׳�6|���}Z>�pC[�&��]l��eX���4e��&N"��3G��_l��l�1�ew�ŕ�*6)P|�}<v��$�|���o�{�Qj^�������gd��+�[��jf�)3��l3}3Ç�f�P���A����u��%�KX�2a�ϊ��q�<�'@�F�l '�����v�Cm(��n>z��;@�fa������O��*�Q�_Ԇ���b�9�:�t��!�1li�Nhl���iy����n��8�L��.m���e@�Q��w�:�eṏ�{�\=F�hO����ؐ���y>lFy �?����L}���/w��wJ-�"_k��7(����U��ʇ=jw����H�ei��J��K�G�+�r�k��X�4%o,Ĳ,�C������χ?��d����
@���9��Y�POSfƖ������;����fTc�ǚ������*��p��,��=i\�s�<u�T�Db(��|0�me�|f}�̒���y��ˣYŸ����i��Z���:SU��S��Z�j�ۜM���X���F�S��B� <xEA�D��\	:��nO��{Z��3"��B��6I�-�>��n�yrS�m���{j$ɬ�F����}���aN�e���I��ƍK��iK��͉�ȭ�P�U֟n�cnG�I�cՏ��X�:�rC�zR��OJ�;G~�N�u��ʞ�2k� )�l4����uT����sQ@W�rI
�T�(�j|F��%*�%�u�a�ٞ�_��"��N�����.1P�EY��:�⊈/O������I��
�9H��0�gW쥫Y��)zH�Љ��}ڴ�+_��82!�T�[8�6�cd���wG���6����D;�#:@�����k� ���T+o�a���o��a��O�~4IՇ�?r�s[p{eFW��1�ִ�1��\��O�4���f��vW&�g��<ұ��/�iJ�IJf4O��B���$�tP׹_~?r�@;k@��zd���R��m�G������c����m;�����f��z��~4�~ǧIuc�A��<��C�/��}�!�O-����޺�|XǤ��AZ'2��VO-n�F�n�b�4��\}Q���Q|j`�"x'�q����6�����i���4?Uq TٽpF���X��2¬�H�j-�v�`���q���n7s%���$��8�/�d��%{go
���='\�Ey�*�?��3��ϛS�_��D��ڶ�� �p��j#v�6�����,�W#}�,%]��s=-2�x��?���E��Ba�9�GH�w�6������A�Wp?P���ߙ��tG��?
����'���WJ��1MwaQa��@�����v�(�����d1.�.k����o%����@�C�g4�X��� �ѫ�����م���ug�̝���=��[m���$�����m���d���t��w{��<�\NJb��o���?��'���J~�dt� �0Ǹ�tg��Y��2��Y�.��9���]�41A{�v{�B )F���K�>9@�v>9mS[�W���#�9�����98/=j�t�����ح%���Tn��m����`Y�hCn@��'�-r���W���B)1?Dd'�F48�,�ë��.&�Až�-=-��o��� 	�YV+i|ˉ��)гL�U~)2�^F�5P���{����~�i\��Z���-*ֱ�W`a��Ie�=�+�n��?����q---����Crr�g�4g�����s�\`Ŀ-E|}��o��s�K�E�0����]@x�4���?a�V��&�3Wϋ����슈l�8���LU���2x���I�M����ډS�[����7иk�iGk��F~C�7 �����(�T0��Ѻט�ǯ��Nu%�=a0��*��O��Nw&+h�s��*X�M��.]���+�T�b ��V����z�u��~MG���'0�Έ9���	��g Nf���l��8�78��
1���y[^����S��˴z�(8��OĻ����a�iz�~�b`���3�@n(s��n8���E҃��p���Xp{)� w!x0!c�Ot���X�.���HZ��z�O&?�t9��O�z��
�Qb���;�����R�.�{R*o�K��AO��-UZ��o��B��Z�%"�~$��E*����K$|�)[�����=_�g9�E�}M�iBN�Q�{�k3��{�����i��Jt�aR��kU��|t5��ܫ%N�}�(>KלS��ٙ| �O^�Kt��w{�a��vq�V!$mz�e�Z��IT��c��:r�}���p�g�0"5�ޒ�R��k�����Q7��׍`��_�Y��sί5�$♜��D��5I���<l��j�k-��sM��5����Z&\��< ��X�
�j5b���,S9�mw�m�3�'���p��j����a��a�H�ޱ��Nu6���]���� ��}z���-��q�T�tL�*}g`���E��zSƯ<���gFѽi��	�v�p�گ�m�i�~��å�e�ɤ��5����/�ފu]�^E�-M%�&��J5X��q0���uKPF����	��-e��l\�HkMN���#�YD��S!�`�Q&UبY~��0���U�����d���W#Cz5(���s���U�e�Z���ׇ�<dUͭ->��U;*b��K�ݍă�s2X�T��x����FG���@-W�nP�b~��a��b�F�E�P�竀�L���ˤ�������&[�2���믬���|�lw��֙/+�j�K�N��]Z+M���Z`"WqEV�Q1e���j�:]��oByѧ�{����hS��ϩ�^pd�6�Ǘ>��$���.1��4����X��j;��ӪK@�9��P�g�g�z)��+�B9����1���Q��M��wS�ٖ��PRԕ������o�'G�0����}���$�Z���W.@�ˬ!+�����|��g%��
�>��1��3��K���,�=b���e˳��M��@�f��	�X�k�`Vnk���[���	�d�ɣz�xXb��ASqS'өB�H�l�Y���3���I�a�{�h�в������]�>f������ �>FdPu�� n�К�W��`	�w�7c�@簎�"��9V��?A��_v.@r�}��vG�4Sn�0郦���5����f��ٰ�GW����~�`j	>�h?&௾b:�����t��O��Wu�/i�S��[E0rsU���F�<���1�"�9�MCKw��|h.�*���c�����6-~�n����3�l�	�wK��;�ꜵ�+�l���1��� ���-+J����6��}>��W��ݪ)J������l��>@u��L'J�_�(s=�E	���]>Ŧ%�>�S0خU>�-eg����@��W����2B~��Ϟ��a5)�d���{®G��˒4o�.z1�d�6��)�G~��jd��&SJs- ���	��R|�D�������o�L'f�����<��Ң�no��[�<������ _nPQøV���%�=�2��Ck^�G�/-͈ͬ��c�R��PUX���OX��e]XX�8Om�Oq�-�8�ٷ�4�-���њ���r!��xQŏ;p����9<�a�ӳc} _�ϡhX���1փ/z+d�����G$M�������p'���'ߗ��9`��|+� |^��D�|���Z1���+1t��g�	���x��s����#��X�!�ݓ-�h��?�"�x�Ne�Y�~����# �>[9�8�/�H��=;r]��i���ŁX�^z�7M�	��x,��G�-�-�.����J2��:%o�ҥge��>�Us��I�v�9��NZ1x��?8�!�%����̽njiaS�-�W�]U�N�z��nA!�mqv��eb��| -��ŚGE�6%I�N����0���O--v�j�!�4����<[�>��aN�;�+��s����@�I�v��O������"����:��1lhci|���.�Mm+�r_Ŵ"�[�-�%_���o"�!x��*�y�+�b�f�x��D��6LE�io-��Z��}v2�2��~o�5Y��"�ӝj��Yft�2ضZ���^��bn=�tp�P�I`�^B�~�4���v!�8�IQ������=@T2�=iς�n��q���^?��+�W����̨�!ӣ�M��e��o$��&��=S�{-'��f�y���m�g�/�����m��f��~Yl��T���&��F9B	f#���`Ii[�Fo���xc�{E�O��K��}�[��k�q���� �}��L8
��'�q]�CI�J�F�K�t'���U+i���:���9%Ă:���%�m��z�nY+��̃Jc�|��[5��F�kV�GNH������=�����hV'�u>P\!��lA�y(d<��2���q��4'�Fb��6����1�p�ݏ{a؏]*Ckr^�8�����Oȸ_���j��I(�6�ݢ���E}wIm�O�	ϴ/��H�����`c@ߕ�C t�m}����A�M�wkF&6�λ9�{���n
�����2�n��e��X0N*�"s����� ��dߥ�����W�j��F���e�.��U�)�;�0zl���A�z_-�&�K!�appcA"1���c���M����yg�� ֻ�'M�����~�}�to���Ā~�Q��N�-I�2 +���]��z���%�.�p#�2փ��Ӿ��3HJh 4���X����x�w޶=��٥��dd��G�.8��P�<l恇����K����j� oM��	���GW7;@�S�*�{��Q���:\6�cUa�̈�Oa���m#R��{#��$=m˞/Rtg�B)�6�9Q����K$$]k�m�3c���0�<��K�T�#�HLlm1&�'�0�g�
��g�_�Y�C�I���v��B���������l&�:�����G~�0/qD�lI��O7��u�L��n/�M����?Z��D��E}���O���J$=�5���rBs��-�
޷�
VS:��˳��a�&M}8��^mE���_Y�n����8p'�!�G�Y�3���i&�G+�y�~�E°����N36�U7����H>K����U;Y���gRU��v��f,+
W�7��ST-P��3��p2O���2���:�OOW���C1�\�V�6�7n'99�����W9`ת���j��:!j?,(�F�H��G�E��F��,@_�we(Ҟf����Bs�.��>��x*��HAZ�m�2�?�>��\(�������?��,OI0���N,w�����0�O�<���^L���J�y�zf�#$��/�;��#�m��[��&����7�Aw�r�t�?|��=�y�w�3dt&��2��K S4W���xD]�m6�yY�44��N���;�$|"
�h�#W ����3��j.��*�f�ړFP��	`����!j�F,}"+I�*ڲ^��5���9vGkfߝ�S�G+����VV�P;ٟ6��_8��`D�oHr<�Q�(žx~���WB�2�:�0e2V ^�D�|M�U�u�]Q�tD���6���zjT��^��~2�>Z��.�z��I����h��J����}~>�Yj������ٽ���l����P2�I��m���6��ٍ�!��U�C���H�Rח9y����O����n���Q�O���Qy3�g�-�vX>S�(��S����ej��h�T+n/�$R��������l����� 4�W�8��.ߠ�bVuDᤩ��ӆ׈|����T�/�;�)��M<F��F���~����qƄ^eĴ����21�3�g��l���[�7ŚR;�1{�HL�����3��mK�llןTW�A[(6n��~���O� �/4ڏάڶL��"�ooUU������H# !ҥ�t�p@��� )�!����<tHw7����<��^}���w��c8�g�5ל�Xk�B]�8�$F]ag�'�������1�i��B	���F��q�����b�2:���>���P��ߥ�w��>��\HW�$�[P���n���u\�HmL��^�=��oD?�Ju�l��&?s��DEX�P�E�[��!.N������c�bL&�����|�n3��S(F(m4�..��X�q�E�K�6����,j�G�(|;���|"���P��SX���_�$�Z�;Fc� ��n�}1|���?�<�rw�v�>����p^	T��V�Cֆ6���io�zct�r�}��DmK�b%c�$6+�yX����%j�=�œ��B�8����HW��a���v����W䥣��9��1�ݦ0R� ڟke�dY�vZ��|�>�u�X���W�@���Mw����L������-�>�	�|�
��Ĕb����2��1*�1�ޘ^+h���%:{�w�aD�J	}��)I��슋{<�}��2\�Q{j���h���)�����>��s��]t�h�Ŧt�I�P�v47p����s_S/�ʊo�d�
�<�D���^�^`f��&��8/r����{X;u�:����(?�4� ax`i��1� 	������[Pj�Y=��-T�~��^�������KP�B�&ǋ�|�E�ͽ�{��a[N�{�b�� 8�n�M˂d��;�t��i׃��N'Ϩ�_�b���6����{�md�t��칄D��^�جt���DC~��.@ ؚ�L��"v�kaq��P=RQ�R�xxD,�����:��z;�V�K�yo�t��"��)��+����QTa������XK�6��J�0�:��N�\��5B{��l3��J��|	C�v0ʙ����\��/R嚈Tu�;w(���Z2��q�8Ċ����<�H�f��B���64�OQNe�y���� Y�N�-�1WNW��$�x֋k��m���#��Qi���|�
&={�'��澨5�smc�&'��:쫇�Z�ߊ��}�X ��5����Ű�\"z�ҧ��x&���v/�zk���)��'�5��񘻸_K��;�ؿ1n���t�u�4��B���G�����zuu<J��_̓��0��`M��.t?pP*��c����h4��S�S��_�o�qL��Ú�1(cj"@i5�_�[�<�v/��3��y�]���=�>�}��x���MX_� <���֨d�Tv��M�k�#&���u;��� �Қp4�a��P�9���	��0���?q9�9�<V�����-�c����-�V-�{
���q�B)������Oo���+�*��������D����gmV�����S�Z�u�r2��|�H�^�&��C�V���E�<!�R޸�����}@~p���[dӵ9q�<r9��.���_�lܾ/��tq(5"aCڻ�p�U�{��Gxa����,)ЦcR�>�NƕGO�L�"-�-r��kw����[֏jD��Ӿz����Ntx�J�I}�D�0�:(�m��}�e��������7�p�`���r����;Z�ˠ�}�]C�>Wz�k|�k��Ưi���^:��Kp0!A�X�}���y[�����Lt��d(�������z���+�K�QJ�+P��K�"��Zw��������FZ�Ɉ�Q97�Ե:g=}�o���J�׳v����
�o`�R��.�+h�����3uH��~�ɏ���O��D��uHQ�7��s�d�;/Э���C/��Mks�u����[1,0��)�7|"����sw��y�:���r�1\��=���Fu�^�,grZ�`溌x���y����I��=��I$U���H���zlgb���.���߲�*�ݠ>�iC���[^�]����*���$Sw�Ͽ�ԭӽP��^�����4ţa���-*>���-���tp���Ð�[�@��.�w}G�i[.Dn��������P_��z��H��MWT�����c+��R������|�癇�1e �KGLkTtH@�i���\xz��2O�<ل�>v뙵�W(�cחBm�$�Ѓ!G��������q]7��%�i@��*~�߳����r:m�c��".Y@չL:�
��͓�5Q���Iw;�/!8��S ��CE���Y�Uv�u���jo\���yD��
�)L��lɌQ1Ab�T>����ȕ�f��9�#�V���\��O!?��l��=O���g23x��1��A'9n�m��`c{|��؇mE�`�<�[��I�Ѵ=taa ��։/o��_��1��S�M9�q|�2\P];�r���ӆ�.�C������m)-��+ق-fn���^o��޼��]��H��k�vK�A�?͂�@�2Sr��ծ�u�4�N��I�:E-r���H�-Ȱͣ]*�B�:_�k��7�.�w1m&�cH�X��|�kB�(�_ 6��F��pa�����o�V��$m��Ao��˂kPd��6"�)�hׅ�ͮ�`�:�$����b%�נ���_�!��bZMNO7'��t1�+j-�:gy�oM�#�69m�cf�tQbZa�,���z𙥓�g>�2C^��\�^�|lШ��~��� �µ�Kr�uӃ��& c���)w����+��f����+~���4qe$SQ�z�d�]U'��e{�hj��Z�~W&޹�;��7a8/v)�*���eɟ1�܀|ۜW�b��Z����mI����bۺ�}��@�-YE�?��I����=t����J`=����c�ʎ���m}��h����(�tV�Z[��unY����A5��OPz�J�\o��a�2�-M��
3-T��"w�0ĳZ�K��"�#(j�)4B*�Q����P�N]֬�����R5������z��R��ͫ>�d�ju�іuK�C��K�(�N�#��p@�I�R]�j0�q�v�}���(A�t[$�Og��s(�|��t
��U���/�{��tz��g1�����c��v&��8߼d.xʘ
mzku_F+�6kڞ�R�z�h��]8֭V�[V�텞�1Qc��!˟P���hi�x�<Q��B\P~Ѵ�5���$v�s�i��D��B�AjױY|_F_O�ժ/z	EۤJ��K�X�84p@h𓙋�g�!>�q8�=�M��ӆ[��OFm`ޝ�
m��P!~��8d�җ*�������	Ͻ���E���̽r���Ӣ�P�^�ܙ��Ud� ���]��<�-��:<��}Ԏ}�Y�#8~/|�s��=Q�_��,�8yner_��	���t#���y��j�W��M�V�l�}�����o-<mWL�3hX�����%��gˮ�lz��J�@T�"�B�.��1ʚm�ԝ?�T�Tu�8,��C�*����/
�z&�V�
�l��hQ��/��l O;u��l8軚�ϩ���,�rW�>U����d⭵:"�NKq;�v�E�/�Í�铁O����r�~�=Z� >�v���E�,հ��ض���zS5��
�sz�{Gi��;.w�b������Z��T�>��5bڱC�����r,���\����ՐY`A�yZ�I�ocݹ�Bc��4Qז>�3xk9|��w�/3|$��w\��G��i���؀r�qﱟ����,f�ȱ�����Ѷ�f�I��b�_$ݮ��ۉ{zI3	�dy䰿rs�<��\Xg%�%��Y����U?�R��������`)�'��UR*��gU�dw����t&u�G�[쏏 �3J��A��,ۃ�q�LN�yq����=z��89�����syz{���C�����aG	���K֊2�bV
^�utQ��>?F�"���w|�=�5��K�母}���$�Z�� Kӻ���Ѥ����a�D��kޟ���]�A��y(DB�	�?�����w_&i����iag#�`�;�8��k$L1�c(Ya������x��Vt^�됥�0��T+n�+Ȕ�u��#_�%j��r��Pc�f�m����K(�cSʹ�R�� +!���(�8�wS�r����k��ڣ�m��$�F��*b�<0� ��=\Q�4����F�:��D��-�O{� ���mx��=�Mt�7,��ah��B���>"�j�8�y�4�Y��� �C�af��^�Se�XR�h�@�3 l}�oV�;�'�3.Ь�.c�O����?��w�S�4pY��%/��|.�	����"n[���3�1O���<v]hb�qw�X����E�6�:a۶][�]���1-���u���?t�ߣϠ
�2,�m!�.�IU�]r�����c���"�p�r�d����,9VH�#���ny��䈠q˕A�l���®+ÃN�����]�~^|�����������[m|�� ���b��=XQ��ϣ��eN�~^�?��F�@���SS�|7��5؀�?<���>���� �ݛv��C~mC���Zt��R_(���_� ���h�A��v��UFScYPqp{���*Ao��9���k��B��/a,�5�$���J0ȏ�Apc_��6�i�%���T�Q���
P��ex��-�x.�]p�ԈS��?|v��0�|��8�7�*,	ց}�z����h�<1� ��/[X�82K^�ղ���e�۴��TsL&e����O~�ہ��~�R�"NT��m������3����3/B�a����Kn����{��f@Y��'[�ϡp�fK!U"Q��~��,q��փG`�Ov�{�"�p �x���K�"+;4,$�����i����tr���_13��/�|��و��at� �`P`FZJ=$e����;ܤ�_��i#DS`wK۷��@���R�ċ���9�0/�j��n��Vr�i����@�y��$�T����ӕ\��u���/7z�=?~A䚐��YiۀH�j�UC,%�U)�tA[�P�%#������s�7a3ywU���ox���U��GL�R���K�A����C�Nx��ԋ�ӏ��,B�L����/�� �=�3���{������v^��Sb�.��<���Nqu9���1]^�| ��k�kk=\�E�ԋ����&�*�b�tL�T:,G��1���?MY���ai��������$�߽k /�[zGŢ��d�O�qN��)|�;d���K� ��2T8ߞ�Y[C�r�,)������0'��,@�2.��Ӛ���ef�g��	��h�K����Z�uYbiS���Q��-�)~������L������g���� �7uN��ЅA�4���Ї��ZUO��{�%;�������`]��|�p%�œh7��L����l? �,��ǫ��|���Sٹ�k���x��<F-itf��xܑ7�]^���}�j��?������B� %o�=��{��se��OJ�~��L-�2�a3�"'�|w�yн�X"���ц�ڟ���?;�1z��}뇋�t|Q}��M��T���6Ÿ~[f��S3�H}�;s�8���7�����3.ΟF.��1M)#-H�4���K��HX	=�y��-a�R�O�e<��y%�������A?��J�=���ɧ\x�,򶓚^Y���vv%��7��j�0r�����D��QE�ui+�8M3I�v�Z�J��-�Wjj�^p5O����W'q�`/X�Y�%[_HU���d'���ru�.F�N�L��p3�2���(���Ĭ'�|;�3*i�BL=��9���O1�x����"�)?m#��;���i�C��$�mx U��k�\?d��Ցٸ�_�4��{��
�����x�B�K�zå����ơ�q矵`������u{��v\!��:[�����z��l���;!�F�mI}�lH�~��wR�h)w����8r,���{������_��n���+79�~lQ��0��x����=Q`;cR�Kj=�ٚ�2�x_�pc��x
�]Ř�	�E�ě�	Ɉ�&����?F��3��7�ỷx
mN ܜ������u�dDBZ<������XnF�я�$�D��&"�����)��h�1wjUs�7p�#<�XW��9��O�h���=v3��M�rU��'hѶ?��B^M�<1'�!+A����LM��ʿ������D��:���{��כ'A�ϯCE���e�
�˿C?����=�#6�?��_G'��gC���[puS7yD:*�^�Pnx�*Nj�K���@�������d�{(���isXF�H_�
ڂ��ɭm��1^�O_�t�{{�{,6�B"����*Q0���=v�����;����l�Kf����[}��=��H��<Q-�ҿ������_��O�i�"˿�8.��A��� w��y�B�ɢ�XTԧ���>�;����䓨
Rg�P/�������ȵxô���e��y�FA'���Y}�2eh���$R~ko[���}�ܦ��՝��s?��F��K�������~94Ew:��������e?w�t�^-K����s�JC'�����q�\�64������&��%ז����âb~^F����>��"$t�wwJ"PB��Vʜ���Z DS}H�Q+�\ �����>2���=8 ��5��E&�C��&�3'y=��w��P��?�s�|,3tQK���<1U��?K
+��kVk��/��AG��,^&�]_�~�c��=*��N�76j����ݞ^ߢ�e���,����<�竣��o9���χ��I"���.�����L���C%ÎZ�;��%c��z��[��B\�"��U��b�=к��7~K�O��S�ǴH�� �t~|�豼����\(0κ9/~j'��x|���64�i����m������U��sټ�W]t�T&�R=�-��Cֿ���Y�@���#�![U5|��̈�T4Ӎ�ܺM�z{lH��1ry!؇�����-6��v]~�J%^�F)u7��۟��XY~�F�gaX�;˩.�Z�>�E��n��z�ݶAb���Z�w�?c����� �5g�>�x�+�K4�;\��4����WQeu6A[3K_䌷��iu��w�>U��R� ����ʓ_Q&�t,�w|R�.D�V�/~/b�b��D�:Q�? ߋ���=�K�9��;�gܲz�wH��U�ɸ�0��=�;8��U�����@�=�0Q�_٦'s%֏��&��3���Ҷvcy�q��5b��.C�V�^N_�RH2��6�v�����g�*'����?a'\���ۆv^����ЧjV���{ 耳��gq,��]�/�)��$-Gee��*���NK4d�T,b�
y\]�w�N�|��^J�l���4	F��ĸ���,^+���x;���Uɟ��r}�}�V�
�qR��"��3w��}��qЕ�ye�t`2�K2F�H;�ΰ;h5���Os�e�m쳦�t��	���D�ذ�\�s�>c�������Bz?cR�jPH�X�����A��C������s[�Y�K|(F��l����o�9}�2y�H.�p���;����cS^}�{�Aq.�d
��fÇ�(`�,���^ر`:��ŏ��J����1�� .5oz��q�����ryt_f�ږ�ڗ��ʍ�Ku	gȨ!�.�r���n�3�J�I����q5�����7W�c5lE؃���i�����.6���ዔ��icC@a��r��S�촵�9��5BJN\�}>%��w$�����y�H�b��*�J���Lp�wH��;<<���6�N���BV�c����V���-�D�͸�y6v���p�-P9�o����6��&�C@�Յ�P]�`����t��.�M��z����2y^��7�80`���&���*�ih-���c�2�0��>!���Sq<q�ْ�
;��₫Fj���>�9��W6���=b�Ǵ����SI9�J�q�����b��F@��R,+=� 1L��x	*��L�� �2�>���rZ8���� 3J&K��'�5��г:~���	r[�E0�Y7���j�R�ݻ���-�0�2��#2;�����:�s6v}��y�W)�ަ��5t�j���o���!�҉S�N�����Ӆ_tm��l������P���K���f��}��Hg�Z���zk�"����A������Ͻ�X��?��ͯ�?�_����T^|0���kh��a��N����°wڐ(��sc���G�,��y�2�p紫)����`*E���X����¥��`�w�A��F�rr�:�J/��S���݆����i����yhK�Z��0�r�kh �b�S�S�HI��-���,O�|��[6T98S�}n�n��k���b���*]�3�I�ui;|�6��������)_�-��6M�AH�o 0�Y~��'���{S�dv�S��kp�(������FAW�v�I~`�W3�L����;j��A��i:/I1����l�6	�w��f�/ȢQT aX�V���	3�x\d�y�-k� 3&W'2ߨ�|bI�;di�P�[,�����]"d�$	��h�UJ{/��y~���ꩆ�����س��;����o����vM�+�B�a�0�'��#�x�iG(�����q�ߞ��UH>��6y�]|���l7����YL<�`��=�-G#ќ���`l�f�h��D))���T��(���u36�����d�vK1,�	E�h�]����b��N��u��U�Um��:�f.e&�T���^�w,﬿ ���SW+��W:@��� hp_`�"�KF��� �0\�$����#������(#�k�V2q�J4e��mG��Z�v �vl�:���Uq�0Ͼ��.~G���@�X�ў�W �>y�&\�L\-��R=��A���4LE�3�u������g�?��`H~A�ԵM{�?UeX(v��i��b㉒�����֑�����J2/V���.��b�Lc?G��:l}��3�f �eV� $��PւF{n�/5���X�6��0����wQ��jt>4�kg���������9��.q��z�v��~,�l��l�_m�,/��^�,��a�����O�e�IfMʲY��NH�E�B��M)�{�	OZ�
��}�OBJi3�));įm�zOo���ELV�t�s`��U&��+�AJ���k������ā�^��l�c���t\��v��b�be���)�gPL!͎�>�(h�*�Lp��S��a���_ SI�dP����G���1T_UU���_յ�G��J��MA) ����(Z�nĀ�@'آ�|��'�4~#��3�����d�Kb��V� ��z�0�+�sa
�z�4�9�{pl}����[/Li1�<���.��t[)�X�@��+ǩ��JG��������g��~�ў�Jo��A�d�I8�s�[°�K\�>�ߠ���dʍ¾����m��覐��v�9��Ӷ�������{D�������(s3v������(�r�7�1O���-�zȜ�B�JjO�l�Uy
p ��RMS5S�%d2 K��I{_��F�	Z�-�HZ	����m�n ��tT��O�LqF{WS���0P�`k���G�K!�:@u� {���#в1�Ҽ�/��H,\`7ܓ�J@i�E�={�����7���LZ�rW��I���''Nmq��&�D�4;#k��"�#%Z��U�	�j�. �H�������y���
��f� ��Je�x6I8�Ɣ
���.j�}&Ќ}�t��Y�A��%���5b��ņy�l����vZe�NW`r��0�旳����8b�ú#j_7lr��`��gi˓�)%�U��OR�!���h��c�Q�Ã�s�Mޗ���;�(�[��^w��y�y�=]w
_��}X���kY��:`���vJ5�n0�i`�s���[����e��Z��{��Q�y}�K�e����hJwI0v��uA��5�Nv��N4[�=�0dYR�σL�ǖ���$���I��T�j��K����E���cYؚ��"�*�L�x����R
�i-���|�7#�QX	�:�\%
���r������L>}�� �v�R��L�]k0����M�[7�D2�I���h=�0�ST\\n��|u�(��a|���ڢF[�h�tŎ5x>�)-��I2�����}��Չ�H���7;���P���.�D]�z�u5'����K��;�SoNkt�{��}��]��N�@I��_�@'q�<��ohy��fTe����x̑�������6�O��6�W!Wu��؆������BJ���z�.=t}#J�V����9DM#���"�$�FNN���R�;$-b~�:�QT�d��������A�a4^LkC�ݣ�Y3{�M�>-I޵�&�͵d7ϛn�_�^�	���rV�����מ�ӻ�rٞu�;i���X���z-����]��i�ДH�`�?��*kH�N�n7K��n(��nh�����7���
Ur�n� E��=��-�ۚ�E�G��x�� �/^�4�����/,���3�ww�VJ��H��w�3\��#=�ewhK�X�@�lfHiP0I��cd����["�0�lͩ�>:���ȶ�T
.�C��C!їi�t\�$zR"�Fd��IZ�b~/�PTܦ���<���`��;�l�`������/��>��^����ٽn�]�n�k��gS�/|U�>�Fk�Be^�A�*�g����W\���##1���J
� ���"�zXW>��[�g�|xm�!�{.����2P�-��x��N��]��9���S��=a�L�{��+FK�"�f�J��{�������S�Wu�i-`��_wl�ϰM�5�<=!�(�QwA��:�V;h�>-5�hΐ,8�2Q��؉�[51��%�hĪ�v��o6���-7KQ�����J�
Jv��F?V�Tw�x��H�P�s��J��-.^���B��.�[K��cJ��,t�%kl�
�[�;q�뉆&�-M�8���ܥ��=�D(�d|��g�j�����y(?�����x�>��"�P_��U�gk��2(?m�D	��D
93K���+N]V�~�����j(i&�`ݢ�5�+2�����������U3�{Q޴[L����<o��� ͱ����Ϡ��!g�^ڇ�n�z��/�|��O�}�L�K�Ɋ��w��e"��܏1�z"��f���[K�6���gj������כH�����W@��H�{{��H��E�+Și��������JK@���UN��*��D��e��7FE��)�&�Z,.��{6���{�4�1�X��C�о��.v)N�:��+Z!q�Mf ��4Z��ߪ�MTX��"��R�B0g�&�u$ ���ƚܠ���p����. ]�u(�ԛZ��I L�m�K�sd$�G1cb��t�#S:ovmE��+˧�/�y@z*d���z彦��IvuWj^w�/7�.���	�U{Yz��{�*0�m��b.OQ�t��Xc����faaf�M&d��oA��t��@N.p�Rj�!�x���o����vgYc���7�5�^�}�S˭#Kγu������➀���f
�eY; ]^�S&~<^��]�ê���|�8�X/��%�TAS6�C�������Qh��W��mF� ���+�>4�R	Ƹ vh`+P0�^{*�|1�����t]��p�,��l�gM~?��<��ʳ5^����������5Eɝ)�-5���;��2L��V�"\��g�����A�G��Fʕ��=�_��]����ʟ]6��Ъd��^�V}����� Ӟ0y�T���gW��,��j�r�����cn�裞�Ν��+�t���ܛ�! �jX�ė-�����d�
���&��9��=�b���%��kx�*$��hfݴF�O{j=�����6�ڪ��F�#�^�f�ȃ�����{����?�w���7�{B'��KWD0�h_�Z���^Bq(���Dđ&�bn˽�c��I��ݓ9Y���R��۰��V۳����������zߣw|�0�fTЮ��pmeo�s�#��/�1�׼-�E�@�6�  #��y;79}��|�:���������j��A�6 z�K�x��k;�ߴ��(�M@L�b�t��B�tݥP�*p^t��[sE�K�s�i�O��1�浼����B7 �qI;����7&�q��E ��3K�������ԓ�Lbg�����C����M������4�?ѹNj�����{_�x�a)7NS?RLgUE�X=�_�w}!���j ��_�'��j�$X�ꊨ�x�^��������Z �Vfd� ˂ZWi�8�4�=�ډQ�M%��7���"\ ӿ8,�L��M�)��V���/� M�:)���@����?�� ����<�w��ZΞ�[<U��n+��G� ��$�T�[�@Q�͐��igOO�։� �0����>NǼ�b��6@;�/7F0]@�~���$*��sy[�.H@})X�ԑ�G9���.��aއc��z1�p��z}�wO�N�J���T�v����F��ܓ���;(�{N<�6yu�~s!3�P`�ڲ �I����a��7�aVk�&d�%e��(�Z��%؂%ik=B �M���ǉPD���ѯ��-��u��B0�e�S���6V��"A1�2<�h�ܭhME�}u�#*�����]�?q0��%;A�Ŝ�.o���K#|�Y��ncw��e�G�"#&WÇb	���m��z���db�İ+l�b��ShB8@�c��n��(�<&3O,�C�1�jQ���������y���h��x��ݴ�B7=ӟ�X�w���$΄��&�/1��m��ZEZY�\͍�2���
!%�1W�)P�(&���N��<�WHM)���䡥揘���j�P<$zm��G����)�>�n@�(B��3�):��q=G=G'=�^Hi�S+T�#�Q4�	)��@���2+y���M��x��$,��2�����m�?�Q�l�v!/ҵ�&�
	����k������/ ���m��SU���%UI)FNV���c�T��TP�>����=���˯_�bV�V=��Qn~��Z�7ƾ��C�%�s:#�Y�4��j��z��R��ǽ�+�'��>&0C�.�g2YP��a���|��Ty�*���k:Cq�UC{8��`]_r`E1�%�V7��\P5��h��٦u!�+����{��ٴ�{�ū!z�bLv'��ׯp.�����_�e��O���Z���J�a�˨Px�ݘ�Q���@E]�ԛ�#����N	� A~�yέYzY��HU3P54���8�T�<{��݊�]����K�&��[�:gF���J��l]x	�����wq�Zy�e^�a�8*7�̝w���阓b�J= MGp?Մq�{�J�.4���~�R�K�m�,X��pX]m� (�_4	�qM�#U����`��L�:��Yl>�~�+yY�Ǉ�������oʒ�kƶ��81��cx$Vy�/�*�������q��6��E:����Y(�k��a{E�Ї
�wZZ�aP�TB���]�ѓ���J��AGĖoj�������@�ž���I�����L/��ʉ��ԉRi�$m�:�V�؂�\���E������pPt����snHW�6#��<�к�ХN�/4�����>�������Y��s)Lum���/&�QV����/�Rl�?Z�]�F���m�fW3�l�~`�9�'��n0�v���ufV�N|�bo��~8�ˈ�#�� E���h��������2�D��q��்}z"��z�U���:0L|���Z���zc��!C��Y����]𢈥��^��w��Vv��%���c�#���%�Ξ��V��Q���|��mp��K�3�q��pH~�dP;�a��!�s�ռ�m�����y��Y���W0�R��0���f!�9Yz$�,�\�u9 ��mL伸8�m�Ծ��|z2�m�y#1ϐ�����4��Z���ʪǘ�s)ot�k�����|���+ D�����ZxV+I�6��ٺ���C�4$��)�ۘ��e}�"]!5x*�����(��������8C+����3#�
Z<��l�宫���/�����pғp���s-@��U���H�U�X��1Ht�;y<�{�늗!Y$�Я{ʞ�u=��(���I���Jtq8�j����H�ۺYG)3&W��&�h�=����N���8�� �Hw12�{t;�L㯚����[�:���m�t��'L���t�.�?���Ս@ŖJfS�6r!��y}L���=0�Z�H� �M`�7��	�K ������ŌPɰ/���p d��~��W=���2P]ě��I�wV)��^V�� nl��U��D�h�������j�k�����;-a�ۣuB�ć�	�l��XAK�)�1����G��F�֔���3;�Ga]\.���I����|���K�M|���#YK�x��P�g��3KsT�a�<-wl��G�����C�E�ʥ���;�Ye	�S�Yam*���ϫ �Io�A�>48�V_}��E��<�2%����s�=l^��-LC�\}�ؒ���L"g��G�Qw�)�}�́m3��4P7���ȁ�P_F�M���;��͟��gH�|:���b�/����`�P�B�����<���XI�ʼ��#���BN�y�"[�W!c���_�3�/)o�����-2���d����3�Nh��J"�lVb�4Qw�YZ�)P��wQN��j�5K)*���B�"n�^�XX�o\4l���n{�g�$�
�ؤC�kb�xh^9����t��l���8��c���Lx�Y���=	w �=�ٮ��LS]L�g�De.��*����GWRm�[�zst���JM�%[�r@��T��y�UB�~����{yS����p������$j{������i�kg]�x�U[�K�_��:������aV"$�m=8����L�?��$N���>��)~V��<o�G'���#,������"
�;�LIJ|dB��=�� 2�.�K���=�G���Z,Ij�)dC�ae����h�
�v�"���<��9�;G�mVa�]%��}�\��n��$��>?�l�cۏ,<����������O��<�K|�`W���>�m�3�G�_Ie'����G�W��^��V�Ψ����I]l^��tM�Ugs.>�}ZC!� ś����/IeU�y��1��>���>U����%�����ْ���|���Ė˨m!��c�[���J^�����	��b�V�u~����w߷��F�A���5�H�Ac�֕1����:��_{w��B	Fp)G�q��-��d��o��!�ٍӃ�(o훜����/(�1��Q$ػ"�t0����oXlͭ���*�_�.���_5�Y��h���P��y�]���O?�d����#~���) ����O��[�Y�wq@���A4<����ώ27�@��d��|p"��#)c�q5�������9|�-��8�C�z�mC��%k��j�|��#FJ/��i�����.�e�d�%}�I�'p�������8 c�NI��=mܪ P S��P���h�Ër��8�o�a��gTk#&�p�9�%�����0�4����\�$<��'x��]8.�f�j�&�I���7������P�
q��ވ�f��  �L��5��u�M�ݢ.��6a���hJ�X(�x��(&�F��Q�>Y�)��C�zSf�]�����z��C�� Yh��t0�N�2�S>Q�o�2Ɩ3�o�V�`R��ŝ���k�>M��=���WpM���F�0u�n|�$4��-v��G0O�XX�+���67cZ�#bp�:hE%��jOT���<"�[]�G+!��p��x���b��=�AB������^N��LdK��L����Ѻ��ܙ��3�����d5�䅛5T���5�u}nFc�<0�j)�����g��F�ʻj�9�nt
(�/k�?P	��f!���/p{Z��@�l��4�'N�qM,IƧڃ���VV����ȶ�~�\0�����v����<|�̄�Aut�L`&�Y�è�JS�}q����Z!�=�.��k��o��a�v���3�w�o%�(-"�vM�B�����O�y� �B˭s�io��i�e��'�q�W�M\�+�.�V�%�.��LYv;nߜ)#{ʿ"%r_�+Idj�M=X����=M��������`j��}5]�=/�����8h�I�h&���E��oX<<��%�Oα�ʽչ� n�w�̈́0P�nS@�c(�`K�J(���_�N>��!N��Y�d]��\Rɀ���Tw�R%�Xq��7�e�P��@D��y�A�����L5O[/p卵� 7U�P.P�Nݒ��t�<U�:)A��h-Ο��m^L|���҆�
%�͓-��$F���no|@.hg��@�:G��4���>�٧ǽ��i������x�T��Y;���q���v��l���t�F��v��Xa���B�b���Cś�F<��Dq8�$`�,AC���"������2\�}��v[_N��z��0{^��!L���ؒ76	�!��m���
�R��a<ũ��}�O�US�fB&�T�>=:n��4ĺl�#@���v�������=<�>_3	:C��t�&������(�%t�S%S1��W������v��RQ8�Z���l�_*�Z#��s��B��-��f ��/�6���㮜w�_.�����E���4[5��*Ԝ�	�{�܏2�3Q�}���M>W�{^I�����+z�q������J	��P����f�?�����^ď��>?�we{I�Q����Q���I���� 	jG�;�,�6z?cx^F�e��J�qK9��4�֫�^s���:���:��Om.4����ɠ���-QI=�nk�-�����/*�2*�m��Ƃw�� �%����!����=xpwww��yo�y�w��#�F��U�j^sUu/Z׎F�
��h��Y�v�'Z/����[����Q��7.��(�o�F��?n��������c�a�*�������mce�Y��6{D��/7�gEI#�Eďi2������^.�Q�bС��G}�D��;~��P�zCyoɹ^�PW" ��+��{d�,k��>��m��!s�˦6Y����Vƥ㥌ǩlXo�%��3���5��}��G�U��st�G�%���8ޜ]����������(���6���j�x��A�j�t��0������A�S�V����&��N8J���RԳ��+\?�W��Y Ồ�%^ K���V��r�m��+_bde���_�\�2��i��by!����Բ�4�����:�����P���@�6���sBEfa���Đ��c���@�ʳ��Q��欪#c�)/��f:��UJ��&%u]������-3�O�J[�Gzz��(�`��h���F	��%� p�G�,�ws��>� ~)���w��hQ�
�΍buX2�7����e�5��E�7�N���N_�?�͚p2�3wwPtn��C�6�r����]Ę���,N��Z\].���շ�	��R�]�
�\�N�kȧz�c����S��nr���|ə�i/VT(&��X�r�o�F��|<nz�afV�s��#�j`X_~�I{N��tXJ~�'�i�כU�G?"(St|??�:n�'��+�w�u��1��}�4�G�vp�~X��O�Sc`a��w�Z��*�}���a+�u��	�J�s/*֢����}��m�_	�ܫ���b%�(�׾��{��)t���1�\�g�>�m�W�n�������8-�����L�ۂ-���ǹ�.���W�;�wv1�kj߬��Z�:/`-�>C�Dmp��͒�����t<��8J�OK����=]]�:t�.��D~�a�r1��������x�'~݂ea-�k� v��)�����{%5�hM��)�P�EdP�ُ1#|�ŉ�߂E�(�z�7�����׭����r�-�3Q�i����L<ޮM���ա�p�����ҡ��E�yL�t2p!}u`�)�Zb�V'�{���Sв�����i�aFd��ѩ�A�ɭ\ճ��7��}�t�Z�Bv���P&�#���2��3Q�,�|̢m6��b�����j��K���s׍b{f����-�	����}+\M�11�q0�{j��;ײ�Q�~��=�O�vS�IQ�I�~Y��y�X�p���S�8���^�A�C�+�D�k���Ā���%bx����n���k;�6�=!��[?�o�;�ƅ{O� We��g��I����>nf����RR�C˘�֛\��tFpLb~8�����5���P��d�)B
��Mҿ��{_,�h�>���,E��\���IŴo����ٓ)J�$�"�~?���yaHV�L�����������*V'W\�و��72�,�se�39��0gpjq�Ƶ�ɨ��.&�\�L#��7�Y�r��{|n�Iptţ�O���XP�
���5��[+������qm�o/9[jGG�hM5��\�-�VO�%��ن4�'Τ�ȁ��ô	1_#N����,D_r����N����$���.ގ��n�}|戀��,ao�C}-��e0�����SozCr�Y-yi�� `��ٽ����#�S�m�u�Z�t}ƨ��)z�c�	&YS*I���'������f��B�~��6�+�m�p�����hjo�_ϊ b����љh�Q��v��n 4wF%�pO��5L&��J���>�x�r -eq�#ɟѲsj�ʮr����ȸ��5�� ;�6O	�6!0a~���k?��Ю�����l�ʼ_��+�����l���g�-"C���;o�QZ}�fcx'?���"�k{��h�t�6fB�}D�k0�#��6�K��4�{�kǪם��E�v�˒3'�}i�P�p�u�X�|�o��Ţ;�(�3x�3_�I�#.z�$���)��o>Y���}X����1�ƘG�r���<��v������JגӬ�5�C˵��Q�3��[��v�x�?7ihV�̟�*�#g��g	w��B�p3?hC�`ևA��U0�1s��ZhO艊_ �y	8��VU���ն�VM��ƑǊ�VuГ�OG�7g\8����u⢜��i^ʖ�%����7c�3�g�A�ye豪�%�o�.��c�} ��7*xeq
U6�(O	�s:��|	8�g&�zS�J=�N��o�L�����66����҂���~�<�n�;:O��<���!�8�����.�������P�L�	��S��`oZ	v.}[�ׯW)yI6��~����Ӧ#�~du�˝���hUl�� �^�������gط���4��=ǵ����3��?�����N8~�5��ũ��n�[�=��T o�	&���Ri/OH��.��v���N_�~%i��X�
p{$ܙ��]��ezn b"ӂ6�J�+w�H����f�`��^��4��i��j��`�/�*�q��H�ԙ>�`T�9/5��m��l`����yY��Si��Q緝�4b��X�#�7���4^�z.��<k��q쿠�M���i��d�|��<�8�'@ԵJ�,��Ym�K���.��c�˸\����)��fE�K�ܺ�He�9��]�䦫(�i֟�,� /�/�ۉ�.��Zl�M�>�Z�w���7G�i�irt	�o�?͸a����o�oOT��o�ܟ��`�KKK�L�-e��*;����^_����M�QU�8�^<��g�}��oW�oײ.ڬ�x�o��n���\����Ѷ=�(��T���[GQ	/�$��heR�#�ɪ./L�SN����8���z�yM����� $�rB�����Y�PI��	F��*��@�Z5�c��Wk3��'��D����0�g�8ӊ���,n<^���=D~.����6�mE}���'�g��zے�sg���m���x�A�ڑٝ��e5mα�sa�����.�T��5��j��X.��
~Qq���2��=�k��,���S"3��auq??~\Wϑ�4'���[\�ź}����3I����@e����6#�x������b@�]Tu	��V���R��mC����vp>��ｾ�H�n�~v���}l~a����>�kHf���k�pPϹ.Ki���J�.�hP�^r�M�2��	Idzr��x���|gw�=6�G8.b,��$?��5�g�vAxF�H�����^|��l�����*O҅����G��-�,�����x���uz/pW��\m��@/W^�E§��ٵ8��Ǻ�`��%$26��z�'���8O%RF!��;���eZ�*���J�8<��q�2_鷌�����?*+R�%�Y��Y�RL��$�ƅi�LW�g�q�JBp�4�n���s*?4��ܑכ�Tێ�9cE��4�Y5>���N��Q2!�3A/��!�)À���d�o����&~�~�"��7Y�`�M�Ȼ�n1;od�V�+�v9�דTf�~9_	?:*�=fK�Ny@J�В�z��m�qs_���	�X�L�˱^)w���iw9=%P�2ee�_�ݯv�|�s�"9=�)�9�ë-�*n�[s�b�ymdG-�!H�/?�1`72�0��a���B�bY�ӻ2��^���F͵�|�@E�s��ڳ~�1D�jvh���oկ̮.��`��ڒ�ҡ�_�'r�v ��w�Ca�1+��{n��B�u��?_����\>m�w��$0n��7�.�� <ū7��8��j�ǭ�u�z�����f��@7괬�>��}�Xn`����_v�]�����F�jn�-\Iύq���̌JZ�T�:��I_�B�c�8֗K��H˿��}v�V��� ��񊽏��Ngx�mB�O{P�y�a���,P2�)���Yj~���i��iN٣�i�������/V�Q��~�uL�ǣ1�|o�O�����vשN��.r���0��zE�۷�B\ԁ~F�F����uA;jp�_��;61�cc[���2���-�K�.m���%� ���#�W�KN�����I[Đ�3�ݫT�Nя����d�d˥<*:���h��s�+�7D��G�]̸�.?�����O�D��D9��	-��2�Q�b9���}d��dk�&Ն�%B��5,P�������'�*'7fi2�GU,��}��'n�MBrXG��m��慄4�Ѣ�`�Lٌ����H�oщ�SA�����T -��U4!����'`޶o���y��U,#�.���a:P�o뿕B��k��H��7�.�r�ы㷽��f#>o����읁.'�~���Ŗi��v��/�o~k��PP�%u�WH��}�xQT�F,�3c��mՠP��:N��v@���N@���9��g/�Y�F!��m�����r����3#	x �4}�:b���jw%���0�掅�׉�p�{��;g~V��m^���@]˶��;�Z��Y?��h-�["�������jȞ����"Or��N��kW嗞������ۆ-�KzF%V*�6}�#�;�1��Y�α0K�+���겔J����-�<WR�8��f�^��L�7�����
)e${�"�5>�	mF�j��5@��Êb�H��~W����f�����B:�bu�^��-��/�e��oa&| �jJ>��U���Jd���y৙o`hZVCy1�����]��̈O�PžIZ�T ����v��~���C��EEح0��"djuX�%�j&�ըBÑ�&S��d��iY��,'@w,�������W�����>nm�"���2�����Z�r�����3�B��~��d웏a�)��o�Y��h�z� Q2����nc��~$X�"��!Ҥ��.l��ۻ:�����Cmn��ٍ�޹�R|$�/�͚��?s���{P{ �}�P\IV������Έ�f�p�3u�p�p �+т~�Q�5 �F_�i�f2Ir0���{�w� ��|�ҧ�(	 �p~%���b�����7�;j��L禷2����7�v�,���X��˚xe��r�QA����?~�;.~�m�����w��ә����j�7�?;y.����j+�`\��fh���i�Z�?-�m/��mǽ[U��jk�W�ƿif�x\{<���3n]/`D��V{n���=Ľm+�����;��={��s�'�gc7xI�t���-���kG���Q�����`	Cj��>����m��;�BG;m��8@b�F{rQ��l�oWr����D�@���>`�5��;�<��vJ?��}�W���dZUz�Z�YK��^_n����v�ly����>����h*o��Sa�!4%���-ˁ��2/��R�yQ���D~ys2����������ׅ�(՟���UK>���-�����ٿ�Q��Y�mr�UV36�zι�)S�]k�g�O�KZ�0�{��������M�?��}Wy���W�/�dp���&M���aVҤ���N��UG�	��[���u��,��<�+�S�Y��7s�jJpq=I�U�j�<�^��VD��W}ĭ�`G�Ƶ�#i}��YoE�L��%~[��?���|<�c̷�C��&�v5�����~h7�Yv�B�+��Ův$�+ӫ5`�&�{�m�������>�w��A0����iQ-J��ϧW/C�{O�����z��=����˦6dn9s,/s4�4��!1:�-s�~�)��)�5{�5N�giw%���������Xn�>(��<�����#�r����8�H�<`�F��,�w�S�:ÍŷZҶ�8/���5�bP*��<��ݭ�	i�P���N�R��jL	�Z�,(�� *�+y����0FGI��B�i|��Y�*�������^,���P��@����ތ�<T����Um��t",���\꫐�xn��)^�O0| y��\{}��D�K��"�A��kk��q��y9iXX�5������T/L�������:�5��|�vg��V�{�\AN$'6��jB�ኬ]m �6s����R
�{v����-݁��*���պ�ӄ,���XMU�l��(.Wr�G��|��9=�ܡr�Q�qְ9��v��M��q��r�P��G����e+W�>~*N�ȹ�("Ɇ9�c�ɼ����w��L��Ⱦ�;�b?�X=�>LÉ��j�<��> �~b�U�뇼.HW{lQD�y+����pA@��T�g��6��F�T�O�/<���R��<��p�"�8�$c����J(t�/����S�,�?_�h���R�M$GM|��C/eϼc�!�DEF.����B�+E����K�v��,��h��W/V�$�}ar��WC\�,u4W>��+y1����,Fыa<��d5D>9	�	�!Rh��"ܣٓ?���դT�]�Z�����;mu��ĩ��aa���O���/�n9c�i��"�_��54�
r���b�<�)�Ӹ��3V�g��-��E���"mX=zQ��a�~���ʏ�M�vp��k�b��nf'�j+�Ȧ��R�.[!H����Gom�_c�;k|���8��#��X�1W\�p�t-��cPq��Q�Z��ԏ���I>����Kn<+:���P���-�@]�2��I)�ǋ��`y�!H����*��[�A,�$5�j�sW�H5�V$SS��x{k��%w��aD�WҴB����/9ٓ��Ѕ��� vg�6�J��h���`��oC� ����^֥�TM��KS��n$YS@���26b�0'8uL}}z��7_�k��?��A�K��O�EhT{�0�/D/4��B�""�G��y'�9�?:y_��jֱ�ᝍ[�����."�e�x���4^p0�͕]}�v���	,�!�`O��Ň���JL�����Yi�F����=۵@��&��j%kǥU�4\�ӽ��n��bK�溑h���U���$���<Y��c��J�e�yl�B�&}���������!/�O�3$P�,K3�9�Ғ���Wh	gmW���I�,Ku����	����-�I�R�ΩԷ��u�.��}�*�ϻ�G��XE�,����V6�6��
J&�uM��Ө��>d�|VY	��&��Q�� �����ɼ��lt��#D-ӳ{6���7��W�v���հ9��L�@J�T�A��#�j'qL=R��AE[︅��b�a��^��M�5�U,J�,t��X�R�.A���s���w���B�(.Y��T��u�=����冘0�~�Mߣf2$h����Nx�2!�Z�wm՛_G��U�1�V�s�ȶ*9��g��(��-�D��&A�t�����Y+8|4����fݓ�Q���b���T��ōh��ȏ�*�?�X��%YQD�$�5��'�s��6|09�
X����ۏ�4�O⥙o]u=�ߦd�ka`�7X���r�/�БYߧuܸ�i�D���O	�'V�S-�_���5vU�HU��.�Y<�k�['�����:'��gY�9�$�ޛ���h�Ξn&�n���e��(�������㎜F:b4�N��_��bV���8-+8�PÙ��Qf��2�'�E�W,x�$��>J�~X�aے�nQR4Õ��,�:�;�����9����R?�K5S5��s�����á��쏶4� S��!��}��>vx�5iC�&۶D�����HPȣ���/&UݵL=�
��ǿ�M:�/������XN6F�FTF�n1��|���*q����(�
1Βy^�
�� �U��z�kk��m�=��~�T5Vf����xKH m�[�������-��#@�/��)�t��{��x�4Y����z��Q#�̈́��\Z��s���|��r`�㵧e�C����A�a*����i���t�q]�F�eʇ�b�����0�@�����ϊ�������Y��O�A.g� ���5d�vGv������Q��k�^`D�K�������1�8��%���@�X�]�#��Dpg�"Þ��uC��<}�ґ%��x'�&P��m�Q�u�������,���8+���O�
Y������8�����2��mP9l�lm�Հm����Y.\�Z$7�Y��� Y�R�f��$�W���+���_	 �E����ƻ�=�kr����>�6M����j�i�����ZZ�*-?ga=gȧ��~�����[Pt��i|AF�}F���C�b|+ݑUIm<᱊] ���@�!�xZ'��~w��I~V�8�7����n4oLޔ<�B�%�LŒ�Z��A�{�4��k�l��IГY
���>ω��m�fX�vA�e_��v#}���i��\h�^�K��N�WX�	C@@B��W�c�H��؃/i�-��9�3/��lY8�e�@aî �'+ȶj��8"�{���O�������!��W`�xE�\�aO(����������0�c�H���@t��d
������4�P�onY�:��MSJ=( ��)�]ٯ|��5)�7�E�
��r��C��js���Hj"�NI_՞z��Pӏ||��k��o���̔ϯXDh]NL��#53�)�X_��៟[}�
��*�7�z�by�¯�2�
}6A���|�=�3���8[k\*�:�G[%��(����s�n8�'�c�|*�RR`��E�{F$�1���j%u+(A�	IT�,�����B��)󈗕��O�v�H`�h8���&�W������?#����l��%� B�"���>�8���aHM�&�C�R�6��-j#
<�'V�/_	�B';����y�W� #�r��� �Qf��TNd ����5'�&���S�6Pf��Q��M��`�L�ǣ���1Q���b��]�Z\���-����wf(�*i�����p2�s��y.4s�#c�aKA��� Hї��!�;I�x��e���u�ە���6D���O�O��9�VwrXܪs�R��A2Ԣ�2U�tȸ̚�%"�%�
��VM�*#B\�W�iˮ��*W��	TS����q�a�y-�Ez�(�~��00�],��D}F8RiXs1�&�]?d`2�T���ȏ�~�&��&�[݁y_ ��+Yh�a��VtX�:k.��<�y�_+���� �ԙG��~N%��� I4�ݜ���J�W��-,}"e�<�����m��,����E�iE�J� ��YVÚ�Vhou�ƓD|K�N�������z|��j*�������Eʘ�Z˱��o�;@���+ *?�X��H����􃖦14���d�׊\����SG2F��MI�lu�θc}��&�����\u��HE�s��;�m{�`#'�����)�1��;уנ��J���_�r���mV3��WJ��
�N�����ٸ��ݚz�?Y����	���Y�W&V��Þu����#��q0Y��t�6٥�m��H�X��1�����i�X�H��y�!>�FSnM�{dߊ��.��F�cv�;\8��<�"4>Z�4��l8=e�@�x��̛�-��_�'��;���F'\>�zg���7�E��{Xx塙 Yjw~����?��|�I��C0�/˕r����R�����Y�4J�OKB��dǵO�(E& ��h帔��Я�͞��Ff��9��2��
%���.��#�b��e�ԉe�^�c�QK�<��g��!��� wl��z�o�:/�����!F�N��]���/�RX���<���������k�,��/���#~;��)��&Ǵn��K�?�gE�l�X������
O$�1�ɔ3���U�[̳������M�r�*���I�a�:���Nv?��rul�7��������'�0�U��G���|�,�-z��[�x�B�����8p������d�ù\����0:�U�/f�Yc���i��qB &�eq��`���B�KC�ND8��i݆�E�ˈL����W�	QK�g�B�}ڻ�$�Y4U*$���w�Z!��מ��[�IX�0G2���U^+�JZ��[��Z��"O/�w0\���5FY-����y����� FVlS�h�����I�2a+v�J�T>[�Y T'�f�������j�1�1�k�D�'<r��Hx�8T�'"�i�H1�;����9���Q�D�.#�!/�O"��D.f�ǟu���a>��8ˆ��`�]�.����|nCB<�����&��_�lվ��gl}m�Ӡ�R��M����-�x _]���G�2vb��nRVJl8e� Y���Z��F�Q��PH��#po�?��^
���Q|S�ϻ��{Zu��њ�{�/(E�%l@"��ρ���uq�>(�or\b{4��lpw�Iۜq�Du��fA�_W���S��U (,��|)�=H�!-��l���O)���|�p1�"�\�~�ՠ��5#�pԇ&�[+��_+���R�z���y���^�y������,q���;OO���t�3A�>s#�ɒ��(�����o	��%�-O��?�2`aX�!%�|�65:H�� +���u�TYL�����џ}�t`��7	q�|(�uD��Eƛg�F��u*���;�����IRy%�����#3���� �&���N��/'Wh��6h>wv�q����dzJ�-g;1f��#+�#�5����¹��@!Jʼ�x@��A�ó���
�}i��`F�������N;<L���y�������wW�$}&��}�<�,���_�x���7⚞�E�Sm7�g��I�� ���r�������=b�e�@C`�r��zP�x��������{}EDӓ���Ә�6L���*�k}�&U3�N+���2�p�n���\&�	���t-՛W��h��Ts2�����K���b�����S�$x0kR�&�QU�LG����qh����J�Cu5S�7̘?CS�k� |(#%%$�ʋ��]5��{��$|B�&�,���o�1�iφ4z���P��}K�J��R26�&T�o��[y���pm7_��������ۘ�I�f
H_C��cE�ٳ�NK��F� C�B�q	B�TC�Ǡ�;h�&��4Xa`N����3_�9b�s	�V ��z���r(w�8���%�A����㘄�<h���Y';#P���=�@��\����r��ݡe�L,]������:�F��]G�n�O��nr�˻�/m�>�v�d@��+�5�ԉ��MC�'�S��5�92�D-b�=������V��p�R*�#�rr�q���?a���t"ȏ9K�):�k������&>F�{�?�+^2H��SR,����a�=(���6{�,7��چH��F,���g	�O"1���u��]cs����}�n�#��F��(��y,�����'�����6���꽎s�_N��釻=�Ο�{{� h�)		i`Sn9�"5�'�ı,��&�K�Y"oU"vbM��s)�:0n�	�%~9Xio�K�L�����H��>7gg�����T[�AM�:�J5T��eP�<����<M"[�K��i:Y�R����UVo�W���g���XU�5�P�����N�ny"���+>i�0��)�G�NS��c����Zh��8�<e bhp:������#S�Y�*����-�+���F�ۊ������$U�$9"CI9�����C�3����:����2�Y��c��e2`�����s�xz�Y��Cy��Q'#�_t��h|�5�G������]��x����f�x/j�n�ˋ��.jXem����=���.I,R�7��&��4�1>t�,O\�l��!�)a����@�&H"�t+�_v��|%Sʕr��A٤ޚԕJ1�`���I:�����P�by���PK@�i�]nF,�[_P`��ǐ9�磵`M�R3>k�K���0V�:�o]��GT �5x�Ș��~�HNJM��v5��w{�����[�,d*s	1�ч��V$cϵ	����y���xu6kz۾CM�F
��J���̺͆�e!`�MnL^P��ƇJ�������40Clh/\�������SD�f�#ƹ3�b�����Jf>||ev:R2e������ ��~�NXR�A ��l]������:�������-���r�%i����}#l4GT����6(�l��BQ#'΢��|��KTMi
wI;xm�^�@~��.d{���^#��5o��n�c���_Y�����r���>�����w��z@NE������{?�e��II��!��.`cs|
a�RJn��1�w�Y�>�Ͳ=��\\���@�X0�j����+d,0%H]��R1�=c���E��yfy���I�^46��$	+4(�P�ۘ�m&���ɗ`k ��#d�)ҭkE�DKy&���;϶t����\��[9m�C��*L���e������'�=5��N�o^>���1�σZ���n��d�\b��G�]�w�,h��l5u��&Nu�ἳ��Bo7����JPN�������M�f��>�'c�˧S� �{ �3T#Ja�ַ��\���bJ%�t�)uQ��M�o5����n���7�j*�kp�l��%,�u�\9��8.�tBf\��O��N0g���Vr� 9�?�ý~w�(Z8C�����T2�~�7�IP����eN�GXDr�Ͼa}��-4<akr��%�T�z��ҍi�}3����{����+##��ʓ�g�3R�&&���#��g;��e���l� �Q?RF�+��w�9a��
N�?y��&i2p�{8�ah?��	vwx�/���p��/b��#O��X�y�-!"�y���&9��H�>�f����k�v[�,(�"�����������7EF��cE���������!��Y�V2���U͈p�.�u�+����"����9�$,׵��)�%�~�q��c5`i�#���/')*L*���29tR�*�������7}LJz����Z�G�&,�ݒ�K�x��7H��H<=�5���1��S x<�""���P��Xo:<����,���~�B�U=�rm�=�'��C��x��au"�Յ�DuE'] &�����AhQ?ݟvz'Ɏ�5�.��x�at<<��N2�e��5$���H�=V(j��rE������7������O^&� H�IK5lu��O*���v>��j�!r�n��uH/%G����E�dOҲ��]��:G'}��o������"[���[�%(,�����?���V�#�s)�� zT7:�u1�5��� >�K	�Q��l����-�i���#ɥ��jc������	����P%��!�F�Y���TRh݅�+�/3��Oغ�jiDS8[�i���_��s�7Wfn���0�N�W6D�M· �g�މm�Tl~� R77�� ����k�hM�\H �,�T��0�n;H`�^=\���}�#}¹� _�ѱ������uh��GZI�؉�o��X| ���#�󧤼����g{+Z��q�����`���C\�H��<����D�}�%�'�~�V�����n/�dvO�Q�Y	����M���a��zڋO�����-�b�������M����,Eǔ���Ž�/���`�)�� �4��|�cc�]��?-�F���WG&�36)��ng�*;��4���\&S����+���gp�rCMK�ÝE���+�v�;a����N����R�,�_�N��q����,�ӆ@�(f�uu�F=b��Yko������L�B�B�co��oʪ:c�
��N�UJ��u̗pk��hr��>S4Դ�΋��!U��=WG�����Y��1$�'Kp�y2�g`�>�U���/5��S�~��fڑ�͉Mp�
>�T�<;}�ҏ�X�����(���w��g�L��]����H�vr-�MI�8�ǹ�A�N�g���� ^+�N>�."��Dr�}ъ:��|�Y�*�?���Q�V
��Gz�@�;�\<�!�$�`�V�a��(���.V�x)��&tK�DA�� ���5�cͳ:k������''�v����3����X��4�u����=!>>܀Ѷπ�hZ/e?.�Oa�4��M&c�4�XʟD�>u��<*�i�}����:= t06�7ҫͨ&�b�0�8��D�f]kD��Xl�(``���
���'�4x�aS9��</^(j����� A/' �?�@���@��VK�ʓ��v��{���ؼ{�'����Ij{�����Ø�+.���x���#夹�D,������>z�O�k���@@�I�Q��-�_b�JA�/�Ϡ�`��PdEJ�e�(��3I&��]Ŏ����T{<����G~��5_{�@'ĢÃ���z�	p��M��SpP�Txˋ�Wk��^�3�����г���Pu��N�mU�z����d嘲m�ۂШ�|.GE�QVh�{���О#	B��������7x�Ǯ���@��~�䉂�|�F���}Q�W������MPd|���E��0����Ĝ���E'߸L�~B�S�@z�f�ס�3���?d�� h���q��[d�@�E����v�Tm��=Y�ǋ�ùz()�����������Z�K5�#y�c������UP�`��=����-r;�&$I�f�@s����Lt*�c�!����/�R�bZ���"�R�Y�����i���E�m�����2" 9W\ ��y?�+�9M!�s�]ΗG�J�.#y�NmNK�~�m{��e����kp�n���QP)�{SuO�_�����[3}�Kp";�B���#.�t�N�a��|��ِ�6��2��NO�d{2upە=�͕��a% �&�;�en`��ԗ�xn�=5�ˊˬ���?�J��u�,ƪ>B䷰�=L'��Q>�=D��$�ƄHP�>[
���Hw'*h�#�G~`�G�"��/�yJ�/u�/$gx�Xrl��/g‬q;�T疂��m���A���kzv�DJ!$.:�������7\B��;�7��ծ_E�����a�Ӂ7�'�0U��)?-�e_���ń�[�{G��2knWcf��=X:�%��W�K��jE��!j�^[Z�O�^��cz���1-�����M�1�������QD�S���':O�4 ]�.Y��c 4�w}E�>�f��=zO.�q{�h9�l�s�$]�ۭ^����ϧ�c�>��.v�⧿J���xO����)Z�u5p�+�ohW�nw*��.��n-X��Y�]D��n���Y�̰���7����H��=��,�o2$^"�aN�!S���R���M;:�1E�Ym�R�$*����6Ɍ�b�1���6VFG5���s���Q����R�o�]S��F�ͩ)��ʿ��w+6C�a��I7��4�`	[�RQ�x⸿3�盹z~1�ڣÏ�X�0|�H֢}o��O�i�ժ(��u��F;P�j"#�2�=@.�?��ć�ū�ˮMrJ����&�����r�����#5�/��j��G*������s�ץ!��#A�u`�t	޶�bAfp���Z"������r�N����XNI[�_B��#��λ'	�E��
Uu�y��Ȯ�su"!�n>�vQ����a����K�r�qwx^3�)�#�XBJj����7�;�~�M楠�K�S\9<%�΍����k,����O߯<���˕0�P8^ � �{�2IĹ =4�<�LSlk����o��.=�9��mr����i�18y�>���c�A2Ի���)j����|z�A���%U���:�N/-�3��B��k-�c���� �7�1�a�A��%2]@{��\�$����W@���`��N_F�R��\�]�ks����)fCqݶ���(J��iD��;dAjAu�3)� �'��a͞�c�D&΀f�7;�-4�{��;�E7����=z武�*M�
�F���K\���]�Qk� �?�����0�|�U\�$�&�8��Fr\��mwNW��++^�OW��W��#��/� ��T7ցB�õk4�3~���<U{g����	;�9��s���T�~]���aj`�H��:ďZR�^��ߵ<#��x���\s�l�1���������"�xT,
B��Zv����ɦ���H�^��ʻ�\Lv&Q<+���|�:���&�Ֆ� \�l<R�[w2N���JK��U˵
e��y���:w�;�7I�h���2>��Uh�bty(}�N�[� ��M��
,Q�$��v��X�KWh1��0�^o�"RV��/c���Kۥ��/f�H���-��.i�+~E�D��×�̯2�xž3%K�٩��*U�k^�|�ɁĊ`�]nE{<�K��r�JHPL��Ί��h�X.Ә�im��g]��U�����j��� me��4yO=��%[X'm2�ًO[R�E��~&;Q�O��_?��_mq���R��'ǲ��Y;>F9���^x"=��yPu`^�R��[D�����H(��x��-�.�-��+𿲱O�?\��=��T�G �m�)�4���?w*�t��̓ޫ���!�D�j|}�20���&�c�qͪ1UȠ�`ǾVkz�l��%m�R��S��BfPY���=�#���v��^�.���-�lT��AK�S#f�$��s�%�;�N�01�:c�ێ��r��+Q�=��%���m�&�nw�奄����Ĩ�� 9����囟{�j�]%��Op���[�Kǉ��H��it7������%�4!�V��vB×�+�oߏ�\4=1�t׋���B����ү{�t�����A^�_�}+�x�R$eś��"�p6��g�hИm,�k&��uҷ\�ty��5�׊\�[�oÜhbW��b��|r�m}eT\��.�	�@p<�K�w���2!A�wH������0��m������ޜo��?Xt����z꩞*�R�VQ�E���/�&3���G�Ƃs�_�X�}g̔�=�Q�4�V��aB���9A�c%ٟ��a����-� _(a�.�J(|�Y�H�i��c7���Q��%��C6M�3�ww<�z�n���� f�]��Z1�+|�n�`:�8I�Uwe�'�/��NL3sѮ6�fu;�~���M�h��7%�1�E�B�6�b����Q��"ͫ��u,@-~�Q�'
(
^�/ȅ ��9���J�B����W�t�`qIg�r�S�&�(oy\�cP7��G-D�W�Er��FM��wqQ:�t��9�Jz�>$�?�����$�ǬEX��ܝ���3=�ҁVg� ������h�!����Vڿ3h��y5�#]鸵��VW�<����E7[���j�8��{�����8+z�����t^�P��Ng�� ��@~e'*n3�w��zlFir��+���d��PòL>0(��m�����qp�k��E��Yb2BQ�ז&�M�X.�"F6E}L�I5u�%������t�*Z�<����-�+&f�lk�F���Or��k9õ���b�}=�)�W0� ,�P�*3(�4��W��U���~k��_�%��D�J��J�c��RR��`��Ϋ�5g.�}l~�}{+��y)}�����gj���l���Ǆ?+bO��	�"�S��8�b��پ[ �ex^�hQZ�S�e�c�,XkBU���'�p�]����~>wD��,��T����E��6^���JD��"�pY�d|2�J�Le-����yO�M���r�f�^g�nS3
LLĢ��W�z��1<dv� t�)k�`0�	jq��wsm��]T��T �?�9P{?�uZ}5��\�z�ʇ���|\_6�D����`����xǯ�ҝ��U��:,�h+��G�E!� ��T�?J~�{�0�,�(Oڌ�U �c���O��T��<|�;@�!��ɦ1�;���z�ܰHe<:8��c����������!�֚r�ߕ�Ո�� �d�O�l|赼ڗH(N�n}��}�o�����7ed��ud��Ќ�^�%a���j�(,WU�����=����**��CYw�$)���~/�&*iy�o�x�r�̛��-1a�7ۏ��=�qAМ�w�C�IG��QH���`t�q컎�L�#]P�^����v�����R%`����w���/.�d�IlB]c�^�!�Lc�R���YW�,DA�(�d�����N�6Ye�<_�;��f?uPN~F������٭yE��2�6_���bZ������m%���H~ ��b��|nC�ZW�܃�|�o������7w���1��@f��=�m�Ê�IbH|�~�9�$<c���;kQv���͖��i�2�S������	�m ���|ma����yN��o\�~�<��q"ա���uf���O�T�5Q��A�¯�GQ�����z��s�g���;��ۋn��Jq:/��qe�ȽYV�N�"���0h�n��m!��<�^؇�X
5pl���[,ϳ^W�Lێp2�nY8a�A�`��'���~�~<O�&xd��t �����_�.::��~�&Ùi�U����s�������|+��|�����NYE(�q���-3�X-^	��=�U��
O�UWA��'A��S&��%�������s��0�1�ҫp��Hg���O����KmukYܮ�$[27_�ƒ��!D��;᳍�/@�_�H�c�o�xfj�Ź�H��v�(�����;l�\��<�)��ƍj��� �����Rogc��:��&2������V��rd���8���7XhE��������ʖ�W�#�{�@�d�n����ÐFoOs��>��6V���X��G;
��ߑ��&ϟ�!�:`>(�wݩM���X�����~ʅ���Xg1=C�7386o`��G��A3��Dp�HM�o�-����c@�8�,C���:����)z�g�$�Jd1"bb��Т�ֹ'�vI�gu�R��g��z�\�� (|AZf��I�!�f�Tx���>�	���/����������e���|�S�"��l��,>O�5��@��4��L؆�O���Q,F��P�W+)8�`?@^�?�*>��H�S7�j��)�����A`z1����`o^���Cޏ5����Pa8�Jy��~-�&7��4�qd��}��+sU�������I+N$�/�_���t��C�-OV�{n
����=c��ETZ�����H;��Ӷi;6�/�u��mO�U�D<V�D���ߝ��n�P�s+7�FB��]��2�7��7&⣯�����n/�wf=�P7��Zg�VGdz8-�0��#q�~����ܐG��9U�Zz�YXI$���*�h𓲓���qCf�ͦ��{�!ǷS�s�5F��7�(l��7ʝ5yݥ�����޶�t:&q9�6)P����2�c;A~?�<��״���6`�/�q�$����i�>�z�!���<�W/$�[a&4����/�%�u��N�����I7K���j6�Ĉ�;ϖ���c��>��W5m�υG��5��ľrJ� ��V�4gQ�ygC{��ǔ�)�j&��Œ��E�ͤ�-��hဪ��k�r�6���!�r����r=Ἂ�m�8��=��ZGA1eW짷�>+���[�,�V.:�=/9J�@T�g摨�Y����=-X��j��~���٪#�O2flg���>��F��_���=�&%�W)_��D�1>�)ɂ�}dB�,&��p�Φ⪨#����"��"�*�ȖPF�(/��ꌝ����C� *'Ϡ����ە[��M(�n���~�'-_~��w5�����nɏ]̈N~Z;���s�I;��i�)�ə54=���iZ�>�94[� Y�gM��������QMj�������+��bQ��\УN#��2WR���V��\v���~��G>,�p�M�F������u�"��N� ���#ȵ�`=s�#���D'Ȱw4�'ثx4���eeo-q�4�X[rxxO8((�T`:�c�);n1>>Rܷ�%��Bm�ݣ��*�K�[����[~�=��X�{����<b��x<�O`��j�/�
~��X�3n8H�r� 㭩x+��[Jꔋrp��^F'_p!�Kkh{ֲ���ܼ��Y�Ї��'�ț[�z��a7v(<t�F��k��+ƴQ��#w����Z������L��2�M�����%7f�#Z�Y9�ۍX���@¶����n�֯eu�!��LY�G�9Q�G�p�Yx����)5�D:J]��I��O�ς��t��ej.0G% )��Z����9.<������6����)�^r|��C���=�I�>&�3��a�����[�<�ځ�|�:��n����|���o0��O�X[��1a5��^�{z�Z���)l s�tJ��
�B�dw� �hH���ݿ�<;#Xn~�����Ł0�����d]9϶!0M��]�U|��`A�c-�eFvCv�S�����+���y�ѧes�/��%e�� �3�#����2��Gzz�ྋ�9�����S�*�;S�AX�V���y����Zsd���=߲��c�K�<�_���,�c������k��Yt���C<�����=w��q�[p�
;X9�����?�ړ���ω�$k�4`�ƻ�{Z�3"yxM"�/�wv���$��ڝڧ�'�U�Ʃ'������b=�V��)�z�)��7q�������v�T����1 ���}w�&��w�[?q���6i�Y���^�0f!�Ԛ����+u�-p�I#_q]�S�R2zү[M��
���ttt�	dS��Ir�+U{���J��2WKU0oƽ��M-����Fk<ū,��6,Rg�0�,xw�������>�2�i�T���~� G\=. cmoCY>��Mx�g��-��F^�����'����nW�w-@[�M��LS	 ���/EuА�ٜ�VT���̸��x��&v���$J艸L�8��k[G��ddW�������?����nie�=��̒�9}����ƌ���o�η��/86�"�-:���,2-�ߋS�����v��xW�����eH% G����ėQ�1[W�l���cN�,�%��֚�As}j�
	�!`D���m�w*��axh�,����ͻ�������T1�U�{�3'��{��^���Ə�؈� i}c&���j?^ח��O&��[�I]�q^�t��u��4�S��'�b|#��9��� ��������D��v��	����ggH�	n٧F���?�l��$2A8������2���Ҽ�������5Y+�^|ƪU&x��}�@B�����9�����+E{��Da��5t��xIu��I����7���ټ�=곗��f߰]�����[���+���?S4T���Ϩ���V�H�f�;�j#��0B8�9$���Zi��U`!�yN�!�@"TÀճ�}lJ��2�kWt��S�N#�;�XM��ž�t��=[��� ��~-e���=t��뻟���9�{����%Tl߆�S��w>*Yl�S"�8�q��=��lQ��Ԃ(��0�u�?aZ'��h���FE�<�D�� L����|Q��ͽ|C�^8BV�v�
�������2w�;��3��Z{-}E;y���V�����v�{�u�q����Z(� 4������9.!#\k@���cI[4����ۗ�gQ�Ry�_��%�/�z~���A�@/88�+�z��i�� ��/�շp%�5����16Ⱦ�5��acZ_���(������z�U6������X ��R^̵�%/���?��oi/K��������7Z�З�䭫Q-o�����	���u��T�<�K�#Z�7�udcN�[	�;�e��� ����ں#�����bM��Q?�m�ܟ�w�3Y<��ZP�I�I�(� ԗ�b�� ���b�3�7�Y�|��$�#d|&ty��/P���c�� A�뻏�m�OY�S��oĳ�v�6"�6��[Bu"���C�*�ّɬ��;��H_|Á�.�m�W����ϼ�N�Ww����Vi��D5}������O�YƖ/%���_m)��ӳ�.�7ZΪ��=# 
�!m��Q�/�AK]k�NRG8�̫vC��V8�:�
䃒���T��XD?H ���0��1����巓��y�T�^$����gy�"t��g�F#�459>r����l}<]��oy&�tW���C>Mzs��<�s��삹��+���T����i������T�����
�{�h�]@����`0w��y��^2��Z�jv1<�<C(�.��E[�e�-��T6^ؙ@���s�L�7�}����}�,�N�<�@Q*(�1|t=����&jtU��;���C�-����]mK?�V��ܞ�D���ez$�z�J꟤�=u�T��'�
����Vk�>�G����6j�q�ׯ���i�PH��M3)=F~���B(���$s n�G �̟d�_�&Z3C�"q	o!��
%�V�_0TPB=���l�pZ�Z-O?�� ���M'-���,h�҈�W:�̵m����eU/XD�Ծ�f.#�	���@�ZU3��»��|����E��uٌ�ܑ/+b��ͳ8l��u@@���:�f:?�э��r�zS�8����{���/G����s�v�'�����Ĭ�ȈF�
�aƇ9�.�c )X�)lW[�����S�Zήaq��\d{4�Ε�ϓ�c%at���7��S��t�zW�~�S*f[����C���|������V���a<����167��fh��v���Z�d�c,&U���uK�k&�L`��,������:�8V�T�g:s6F(,��!BZZ���2R@Z�<�B-Ɖ\n@�#^!�?@��<�s}�k{��G�N�P�[a�Y���L��bx.117��$~��J�Q�L-����zD�c.P���{oyMn�'q�?���Z�� 0���Ů��G���ϳN�g?DJM���$�`d����h��G����,©B�rlǱ�Ă���E�!f�שbH�<{��h� ?�Bw?��}�si�i���鬯p@���T��"h��KB�<�sh�[�o�,�%0�
3r[�U��";�
7��_����;+�-�z7�Q���3��n�kP{#J_w����b#76<Ù���"���� ~��Z�����*5[����|̙J��{�+��*���)Z(P1�;'4�NS�o%bW���~)ob�­���=���0tk.�A��c�/�Ҟ�ONr��?�<��������|��Ởh8t~��y����ƍ0�0��`�o]��i����ueP2;U�������)m�w���ּ�&��MMsVg�y�MK���G$7����� �)O.R-�7[w�CH��x<:�C��jI�U��JY������z�����-]���!$5��o%
�idc���Ncn�;��V0rS�GʻŦ��S}��AH�~U����Y���Y�r����c�X$o|<�(���\*��v�;'�@���c���ί�y����F1]�f=5Qʖ5�?M��s����D6�G_���Q��ݚ��Փ�76�� L�6��K���Z(���9�һSA�5�}�ɏ��I�#nF�x�9����gn᣶���W�(�p���b���F���p��K��R��Jc��'��a�Hq�"S��g�{�f��c��%���6����N�^Sϸ~c|�R��m�<�2��D~ÎCG)ɫ�CmH��;x�7�>�]��Y��[c,�4�/�35d�_�#P�8<�Ό��^C4.�|��� V~n�(>S�W'>95V=6�ɟٸ���%"l��e/�N�#E|�q[6�y�,xz�6D�&J�N��9�-��ȃ�r��_���:�d�%������p���g�jQft�Z�@�V����ߑ�#�6$�`OX��}��Z�,��#�铭]j���5�;$L����!2��1�EI�
��|�{T�w��%FQl�)�ۢ�|6��冊C�|�T3y�5�êTM��������C���r�V�7 �?��t<�m�6�l���,�S��T �jվ�݁&}A�<������N���	��W��O/�غ$�o�,�W(ϞJ�m�
�#��Tc�?kW˲21}P{��:������[�Z�ْ�dy�"�P�Gq�����W���<�|��,2�ng�j����Ԕ��h#È�L􈣞�#$��
[��^m�>Qi_�d�J��:Y�� �5��#����5�g@1���Im��n�'0/G�6�6��T�I�'oT�Es�iBl���s�������4�iL@-��"e'��"�])�.�����fmU0ޡ'T�ٷ������j�x�������xd��MSj$Û�;D��`�l�IiTY�DѬ��7�WzI�ZZڈv�m5���3�Ao�H��%&m.��+�>�>e�h�!.�"eG0e��3E��cD_���u�䃓���iG�-���e�ע��A?�{{�ISBo����m�fU��6��[Mi�>�`�o�&[A, �ʇ��x:��z^z̹�.S�S�S)ڍ�ݓ���j���ۘ4��&L��K*��\7����nI��vM���x5��v��c�Z; �M�SA�ޮ��_��S�jr��k�;]�F�o
k�]��_�^�j����*t[d�.��DU{�\�z�1�ӂ�ZB ���
���^ǹw0p�څf�*6BEa����g�����OW\t!����Ǘ�/R{��=��(8����=S���7PN��E!n�a{4����Jl�a��?2/צ����u�H�x�?"�rlzҷ7�p�ld�(�җ� �ﺁ��
� dFp[N#	�W�
6(�F9Ö�+��ht ���[S.$���I���)�(��x�*(_]�����f4�h�Ǽ��K�#�)��5�ll)-֐01E�я~�x�2^��=ON����`�m�1��� ��Hp�-'\0��C��]J������Ca�Y�:�ɷ��@�Ab�ꯏ @�m�q�1Ϣt����JE��FW8n�/�>*�ީ��k��dy��1�;�m0YX�$��>�h\��侏����W��%����-lxϼZ������Ĕ��XYE���6�i���w�O9J>��}�f_]�FP�`Vu�5�b	�5]CDkg��1U����>��D�@��Փ����Uj�d� (QU�Þ���V�⠟��1�s33�r
 �5�^��J�]��B�񏹵��TN�o�H3�w�'�>��~X��F&L�T�0&Azʬ�+T��Bo�$!/��F5�k~24M��;P���B�X�ēb�� ��9$�6(;�}���/$l����K*�o{���E9KΙ����|/KFSBbrr��]��*E�i"8Mg��tSC�;+	���t����1��F�U�^������̇I,=��Z���j#m����T��g�2ebʡ�#�~ˍA��C��K�O�S���[��m��<6H.s�Wb�>���	�~�>��E�7Vl��/*�e<|Z훦�������-�8Q�W��5�r�_*e��8Sa�|8Yˠ2�c�rޟ�.����f�)�c����^Z(�IU���Sꗻ�C�	����apa+�ll\`\���9�Ĝʦ�q�'VJt��9���=���տv�W[z�a�m]��6}�^�˿�aN��P��e ;�5:�o�Zw�w�.]n�T�\Z�q<E>�x���k�@��3���P+������Mp�[K��Eg�x`�=�X��Eȏ�Ko�U����ؔ����n?ۋo-���r��-m��ߟ:
x���n�J��1�qqkRc\���;9�[{=�kw�\h�l��j1j�~-�_9.�E"�3.��[��n��n��`g�TX]h?�%~j�?�zVб�L��_� ���̬��J����{�~���=!���:ۺ0v�U閺���I��ڍ���1���nsa�->E��?��㫩�ٛK��E�_rJV���f[��ޏ��&O�^�Ɩz���)����i�p���&�$th?�/5\�xK%D����>���S����|+���c�M݃��$+/���j��|�N-ՎY*���h��t���tn{f�ux}��	�Vn<�+}�rf�0�2,�ꊮ������{ё�s�e�|2(s'p�rҬ��w!{#/k��	�eդɳs�ݍw���S�q�b��|���3�V�R��U�t�p����G� ��XdG����/lI�]/�׈eك6�J�x�r��	�����/��j��Z��d�J����v��f�R,G��WSN��<E��C�Ƚ�{���i/HɷOk�!��U0^E��6%�oӊh&����0~P-���cǐ�uW�ש���o�t��"�N�3w�G�%
G �{���K^P)���U���j�k�0j�1��|^�ڈ�-�_���V�e�Ε�M��<��.g�!݇�D�b��x����Q��m�ZQc��[_{֦z�U�ʿ5ldR��0,<?��쎵{�q8F6���]2�am7
ޢ�xW�q������<���Fu���I��ڗ�����CN���[\��� ��{��؆v
��W�U��l��y�j�g�r�HwXCj\����"����uS��!Hc/����B:k8!�֧B��x��p&���QF�����}���E���L.�x��ir)� +��ᾯoX�\k��k��=�A�FZ�Z����ٯ'��k��i�z���Y�k���@	�'{�F޷�����'�V�RN�d/<O��3EҧŽkK��	�a^��9�EQ�}����ʢ'w^�=�/��q�$��[�����B���\ؾo���Nu�(.�^.�н�����\vy��6�����֧�rv��e(�,E��T�4b���W��%o!�<ﲎ�_c+L�d�j��'ҵo�!+�ff��ETp?����mυQ�b�R��-��{yb���B�7������I���K/�h~5�Wiv^^����sf��"�[����K�ם����p1�76�N�����9*S�����Af+�X�`8E�"��V*�-y�R���^J��������������!��z�ڶ�8�aF�5;<rX��$�.j��m�e���jw�Mi�+bO��E�#��k�vM��^d郾E�[���ݔ�~������Q�F\�:��vϛ�qǼD(�੩���������y�5!��p�x���Vc��*E����L�y�C����=V����E�������a���x�k���[��F�$E�I��d���|��+���{�b-��{?t���!:J��g@����l�i7�j�v+�����I(�������ZN-��@�k3b�u2<��չ�}�@
�K+���}��7țE���Gܐ���q^����5]��t�^����'N_xAN6��<':��DI�ْ�D��!0�����Pe��B�[�W]+��)P��^�u���,A����ޙZ����G)f�=�w	2�ȗw߈�W���LF�N<��QƓ�lZ��?Si�p:�C� ;`U?+�H�O!�>�.�R���}�P�ݱ��~�'S��B��&��HT�v^R�(�F��9��!���z�e5�*�_���DtuJ����z<���s�UK�W��F=�zB��8�1�_`;_��my�h�'��+5ι�ޖT�2�g�ms�q�F&$_h���O����_ך��?�.U~���u@׿k`^�?���.\��`O��w�}�az��x�U��� �[��lU9�z���뎸��\7���{�9GyQ��x֟,�%X�q��[���H��o�|AQ[���;h�ߥ���s�3p�^��Q%��&��?�S�)��&a��r-��!&���IK��8�LeY����6ԉw.�jZ��jͥ4>kx���mȻ;����]��?��u:� i�ᖜ�v0S8S���t�F��fƺ�p�l�4�w�	�G� z�:�gm��<��j��z��b�r5�r��^v����x8
Ц�j��������הy%���л�e����4�j��w����A��[�lC�'ds��S��x$���qKxώ��R��.�0��ҹv���)�Ia]+�ݩt��Y�uO�L�����x8H�_V�xk�zfxR�%FI{v�_��&�i9+Q���į񔳲F��~� @B2�)/?֮X�b���,M�NQ��,Lu��e�%M)t�.э���w�n�*D�M�����قc�I�E��"psH+�i_PVVVE�8e�G�� w^�lry*/(Ǌ����Иh����Jn�I�J[>��l���+5��?���Ttu��T��ȥ/�	y�d"���9 ��X�h�h��2ڗ�Ʀo�e
Ξ�k�y+�5w%1���_���"� �-4�n��,���bd�o�q���v���9��WH�g���JIwz�޵Cl���r�����O��(�5W^��u�s��Ǚ9P�j����.M���8��6���������0�G��OEo�-�iA��I��n_��n�v��8w#HD��J5���h�.`=�ߦ��0�Ey���y�����2���Ԃ���fm�����L�>��lw�5Ħ��U���DZ�|�>E)���ջ�/�� �����q��S�K'x����E��Y�F�ۀ-lϧ����J35��O?}�~���Z>�p�Dl���[����UД6��Ǭ,i�QQ���;;�Aϐ���A�X�bm㢎��(m�D	`ޮn��Y�2��vx�W�"��6 {��L{GJ��_�{M���5���n�|�z�ͧ�Փ{��7ç^��!m��)|T7���ƌO7�����t.�g�鷊�fcPw��ysӸ�2?%>��һ>9�^�=��r���f�0�9���~֏���1��Dc�'HHxw�Z�ļ��ǥ&C�sSE5�&V{6�t�Stz,e�aa�)Pgki�jX�W<(�3� [�	��{�TLƱ���"t#����,�Ȯ�zV�{n�Y�lTU�WW���3���⩜����:�/��O��B$x�#�\�{&�2��6�e)����8���@�~=�H�ކ��zo�5�����c�Ґ����)�8� ?^�AF��wB�C�G�HH�;.`�+��Y�����L �m�%���U�&�53EL`�1��	=��p_<n?�A���J��7/���rE����ii�q��\h�'G�Ͳ�1��Z��u��[

`lk5��k}�����Euy�$�8-EZ.��~�K">�bt�JGf9��=�`�ǋ�*��c���n%Ā���F�}�^8���K�*����P����,������l�D[���EM�?��B�ڼb#ldڂ�.g��2��a��~	��w,(�XH"OH;��"�VN�"bL��K����0B������oE�I�f�B�Q���c?�.��_��c�/?)�}]� ߼�+^��z��	�H�x�M�@(H�y 7�pZ�Ԭ�0�FO-�<����5������_sK�^ϭn~�����>�Z�ȩշ�M�.,:����,�t��Z�ٴהP���MBf�:��]�����[��+�Z�!(z������W��Ojl�C�� ��3�٦Z����ðA�dJ�wm�қ�t��ץ�������p�s�Vd�IzȒ;�����PR,$�:��s^�L.E_�G������p�`_.n�B�J�7��V�ř�'wj)�`_�^QR�����Gg��Q(Sίj�b
W�D����9z$��kui�Cb}Oo��I�g�W2~�u1�6C:�E3Bj� �$|�1 ���l����9oٖ�m�p��a��:`��1ۅsYM��X�w �"@ދ�\�}��.�扏 }��0ac?n����9�{(D�͠�Ak�5�U5`#��D�kV�Y�s��צ�v��������h�4�F�F�ɩ��	�jTs� ����D��,���$Z��H
�ϵ�>m���W�(��ok~�Q�[�VՓ���}���'rC�5�w�ۚ��93@3Y<��B:��L˯최#�� �:BU�W{	Ҟb�I_�JXx��]��QL�u�]s��!��ł�xDtohС��	�:_�j�R1���c낇e�.H�-�jGn'<�P�)����#��_7}��h�%�lY9���_��+v�]���#$����	V�2���r�3��=F
��l_��,$�p����ža��Q?�J~r��O9S�Ap@����)ߝ}��KE�?��.��q�-.�Rr�Fc�x�oiI�d9F4�6	2�ݘ��vw+�տ��ũ@H�}S0@_+\�7g�ȕ�MOێ�`_O�$Z��R�++�i�0,��ظ� 5K6��v��3�ޜI���qb � r�.�����?�l�iU�;���u��������F�ț 5�Sjw]\`%�����8�|�����>9=�^�^��O���+=_+zuqc�ɑ3���/i@�N�7'0�vf�y}�d���NOZ�¼~���St�4S��?����Ts����4��l�PH�$�u��t�	pP� ��~ј��s���nh7�����*x+���j�AO�5�jŔ��1�w��o�cڟi�84��E�ع*9��;��c$H���)��Aj|~� (j�X�Z�yr���.m���ZJ,��a{8���Aff/^	2-�s�]�ԶS����/��6������ &��pY�� 46Y��w��D�*̉�	�K+a��A��v�E��VG6���I�(�NO���$���R�<� ů(��x.'�>�Ep���}���B�dW�!b�7�d)�4���T��.Z�����Mo�dTO���K>�;�a��g_d�|�ۺr�U�]���M.�R.B�C1v������TG�A�/hC}�bm���Oߖ��F��"1�+�
�u��"�M0K���6��T�:�9ٗ(b�
kfI�I���U3�^�.!�6Y]���E�)�"g�6���WЯ�E�lf7�n�^��Y����?�$�@��Bz%b�W��	�\(�e�k&��HL�|t��J���Dr5�}Q2��{rS:95Q ��2`��T��(ø蛀���J��c{w���XDJ&�Z��� MM�˾��&��Md��D/�պ�����|j!{��r��	"�0���,�g~�a��[���zx߾�|?��ئ��N���ϒ�iu����gb�V$�����,O��c�ɍ��)����+��_c�*!$;bc�5H,���J��L�w7��~��y��1�@=���܁<����^��[����c�>˘.��sB�^4��\�먌��CZt]݁�����	�zE�\D����n����s��̢� Ӯ�թ��_��8����� ֯��X�_��4���i�1{�s�g��Y��i����}�1D�B0����.·��g�E�B�lJ��a�2y�i���r�Pl�0].mӚ���;e���dT�Ǐ�Z���Il�`���Wߙ&�J���5`�	+��@M�Ҩ7��P��t̿_��A��
�;9M\�zO����lO��[#�٦L�����i�� ��ل�h(Vy������ ʾ�3�s�1ً�}Ϗ���S�_J�x�oo�2_J�Jdrr�[�VU��(i
��Y1�n�!=:-�X2F�G�:E<Ѫz��sV.aJ#	OcVǖ)�#�,��U~�v�����&k
cW��F�x@��t�eg���1��Z9�ze����מ�%
��K���i�z��T~����w�ȇ1��5H�㽄��3{l�$�.i�y��Q�ZA�댤�"�0K˃�>G���__�0�eoG"ٔ*|���bIX���Iؠ0��s��oA�ڻ֢�k��y��X��Y����",��;m��Y�"[����"���N#��1����<�v��}NH�9�-�_��Ύ"ɦp;�b��r�)�۵�T�N������m��dl'�eb�����U�|�]4C���M��.�l# �ժ�q��dv�$-.j����%�cQ� jr�ݵZ����z�a	���i7��l�'�ͯ�9w�9�M^e�3=�Ԃ0;[N�)��{�������򌲜��Aҕj�m����u���W�I��R��J�=�j'�t�����<�R��^�w�2u�A��Z�P�A��g�Њ^}y)�r'9s��.l��B4'��Ѱ�1�g&U��J����H]U��]o��1��M�2��.���?al���B��%mӡ��b��Q�����+AC��Ȋ��9L�8�:9e��r�!�C|G�p9���m�^�޿7�]�v �v�t�z�VN����E�� Z�KEJ1������4�|���T�G�2�,	6�ʶ�뎩z�M�`%����wt�JwBN��������C�Yśs�q9+$	ߨ�2�ӮSU�i��{� gg�̩F�]b�C�^^L����3�J����%�Mp�מ17E�#Љ|�j�j&�����[��W�a�Xے<�s.�. _�zB^+p��{g�Mˋ�L���X*�����v�WU�����;l��J��<Bu� �AvgW\������T�|L��8��n�=�n�.�H�IPzp�l#��U�TEB���9��z\��I�V���ow���k���WUU���r\[}5����T�!2V4��ˌ��n `δ:Eo���=�vVB&a���.c5��]���ۖ8�*RVψ�
��nLiJ�/#NUu��Sy�;E���dWY����z+5�uig)�x�R��;*��EZ�� �=�yՕV��d$�u͋��n��RˁY5���:��ye�#b|G��ޕ��Z��Snk���;��
"Zl�%��n/O��1�@�{�? ^��lF��-(G��0lFB��k���d������t2$���/2�E;�E]�ꖩ�6+3ص�fG�uq���;M���%k⒌�I��l��[LG(�2ߗ�5�� PK   `��X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   `��X���  �  /   images/dffc241e-8a0d-4217-bd54-7504444465dd.png��PNG

   IHDR   d   �   6ke   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]x�U�~g&�$@
	�PBK I(A��t,��
���eU,�k[uw�u�W*�`�w�7C �@%��:��=��If&3I0�0�9>W��/����v����°��������2�0܅����Ý��W_Ƴ,f9��2�\<tqdbY²��,K4��Ύv�K,ϳ�X}�&��,sY�࡚�؅),+�>�'4O��G��dy�I߱Le����,�X�8����Q�Ph���= "R/���za�7�&Z~P��PU$��/�O�,������|`�n�t�������� R-/��zb�_�h�o2�~�>��I�Fk�
:UG�y��fr�ZeH������������Pu���7`x�������,�X�����2�Fk0|X��CՑp�5�rfVQkl$ChKW��k��0�|��mB/�\UGb�byQ���=/�Yް�#GnohA�tV��ʸ����Ք�͵��I�g�H��,=���Y`(�l&{��qh����@x�b���Y��y,�� U�t�g�3ՎD=�Ƀ^�[�7# nF@܌<��y q3� �f�������7#瀔�	�t:�S�%��x�ܭ�}�&:��[P����{�2 찏��;�Fx��0��� jBޜ`I�9�hD��Mɩ�*�ʒb,+�&=�E��c�݌<�8��ؙ:R{Nѫ�~���I�P�T�p3_� �����+(Ҍz5�x���+�1��(�'/FX�M7VO����(6��Fp����6��:�X��C�����I�p��w9(�a��%�vwf\sU�L g�ƺ��GydLB�����">ə�УM\ѱm�'��}�;�O�X�7�SPPT���uf��q'��D]�c���E��;�C�Q��JƱS�x���=��|��4�8~|�������0w�N|�i��v�㡑�0�G��yS����_�̡��|���۱`�/HN9B�Q�ƽ�Y�x���N���"�ܟ��w�̒���i`�;v0-�36=�F(�U$A^>g�ZJ%/)���	)U��Y�/��_v�#�Y0���IC��F���3�ߦ��f�$M������{Y���䣘ԯ|}*���`?�/��8{�pV�m4lR�#��Y��4@8a���'��:"�K��Â��`�z���a��=1aP?�3zgdb����z�O�=\I�aC�g�!>=�"+��cF�Î�hlLJU���vG����*�}�֝�.��+~BN^>ڶíW�t�2�0Z�)-E�L,��:_P��o�I��R�������2v{j�b�=��p�>1jn��]-�D5���^&C϶-���k�s.-�()v�DP�b�2�M���'���bad�K���c�>��	��w�bϷj@8K(!h̼�p{U$jL�ӎ�V�)��e�R2�)�c�#���
�ye��e�@����]�'S�⮡m�@[��������@t8I���Y�:8F:����&�eF�)���M��#��=�R��+	¯8�}J}N8�ıw8-�\MU��J�v:�͂��>��C����1p��uz�&]���`X�Y�&x���x|��ŷVM�^�������NoU/s�q�sШx5Brf6;�v�A�1���۝M���wmB��*5�rB�&N{�c<��Wj�j#ߝ+(����ց�U�TAI	^]�	[�������0u`o>Z��xӞm=|�^�&�� ���Sc�Ftxh�c:���cCU�lI�����X%Ns��*A��U�d���g���Թ=��~�:�N��J1o�.�QB�5��9��[����֮r��S1��UHI:��h󙰈p<7e"�����\5���4`��Y�疟�BAqI��Oݐ�I���ʃ2�+}�5s8Ƙvm��iHL;�َJ���M�P4�kD��̓z�!d��H��k�H����]	�9��Hڽc�ګ�jH���パ1ј�a�Ũf�5Pb�Q�%q�[��1�0Z���$/��j�H˾�0B'�$&�ge*���Q*R���ܵ|�u�_J�1�O�2�)Y�ۺz����<=�8��9�w��S*l#�mk�|�-��w�Pk��@(/ˮ�R3(�l�~H}�P��Ġ�v�m����Lp�[���`�XѠ�DS�z�O�_ޘ���^#u�7�5hA�t�Hʥ8!=q���wy�h�c��]6��z��u�PŃ�.]�y��\�H]�#h䣂�'Q����z'%��j���S�ơ�Ұ�g�'�*�Y�u�P|�����8K�����+�1�Ǖ�3.�IH�������Jߊ�[Du!�@�i1�ըH������F���SD��hI�����w܌����]/�)z�NL�C��������b{-;ԕ�ď�F}2mI\dD�� ����Lݸ��N�-\	H�em@љ�.��.�����6a��җ�U��6���c�"���
�q�]�lMo��~H��35�ڬmp��W������!��wf�ۊ���(=����6�����9,A�$����^�ڹ!M���b���qXv	e���O�F�
s�����:��M)�e��e&%��P�y7��V"[��*u��+AaRF�����	'��dZ�JM���s`ſ���/f���])G0}֧�Τy24.YgsQ ����ju�\l'!"]Z�i����| �i2��>0�n��Sg5O��w�W���ű$�C��3���hᗄ$�B����>ؼ?�چ��jw/�h� 2����5��/�1P�94��P�6Dd���}Վ�,9��ضK�%��s�t�(}$Rh-�Wm��w}��l�O��NWoųӽ3�w뤼,C=yY"����o��R�]�eY������:8�c!�p��� �Ux�3O�+��6���)uA��0�&���d{M�9 �xة�:�h����R� v��o.��Q|}0�[T�hU&ǀș�.ڠ�����f��¸�n�P��C	�%8�O�D=T��Ԩ�����0���B�_�{��(�InG�W�dn�2��s�2�.��#DpCL��X��߼e���7%�������1����Z���4����C"�	�?76�(@~�������7# nF@܌<��y q3� �f����) ��S;r�qU��L��=һ�.��z��7�܅��*,-�KK֫�jS�؟*'�uq�W�C	�s��j������ ���!���r3� �f��ͨa"�:[V��.G�$i��ʫk��5n���X:&-�����>s���r�=��\xh3�2�J��)�hl��R�%�aB&�m��~z|��p�X���7�a9��䭯&x��)X�;�S)�������Kr�H����_o�9+�a��_��<3�F�0�/I�J�7�R��E0~�'_,R��n܂ןx a������x�A���rDn=����--Ųm�1�W��%r����;�#΍M��E�2"�`�x]�4H@J��%��G�ޫҹ�Y��� ,ٺ��.P%mK<���,~�_Il�p���;�!�"�n����H?uZ1�� �	Bc�F�v���$@ٕ9?��Сk��f-�/-���$ &����� 3�_�+/�2�JҘbԭ���g �}$�z�n�Q_|�jr��{$�eDF�;n�n$v}����pǫ3�G#��T����"-;a���]dy=�D��s�Ԕ& �2�t����	�_~G��{z�x��a�P"ʳ2P�����tu�zc
r�0��>�۟��|��*�I��� 1�[
a|����PDճeO<b���;b}�����G�SG\�O���LA���hD������ �"%͒�&zP���e���%$6�=��X�/��Gye�lڂ��y�dϤA"I�۷�,j�j	Z����X"9J,)1h�;0���t�����x�o�����z�.�v�{b��K�:�U�IRZ�q��<7o��ѮU�eW��W�ñ��xU�uj�޴��� ���ٹ_�&��kC-Z֦�N�} !�t��*Gչ��A��"��J�a�0m���=g�:���(ϭK����?+��1'�����Ø��[�U�a#zw����<R�� �O��=�hw��P(v��u�O��q9c�G'�QI�l�^��*'�Ty�L�l�\و#�(���V3Yޔ�}0���/'~�غ�ϛ?������:�3���v�Txe1����n�A����Od�R׽�x�!�|�I��?�I�������n��#H<z�b�j����LRK墂|}�^�F��t[�Ȭ�Y�2���9P1����c|F�	 *�U���RR��V����=�).�R��4
��?�$�	���9��rx�6H�[Z��Lv��N⃅��ѿW�����T����K����M�۸+w�٬����Y��d���#��/TxZ�LQ��&+5�6˩���m�=�l�eI���ڥ�t������O>�~����a��L���djD�`�>�"��x�%��()�jSIU�93T�+�id�P�Q$w�RzS3�>���{\��ݥ6�Μ�Wu�mxj�|[�.�ը;PU~�����I?#BC��/6e{}��%Kv�D�zK��K;(+��_zG]�h�!�b�&�r����	cɼ��#	�����a����Q7�	hr+�F�Y[X�2��Ոn�Ryf�D�z��Y�@�!���m�wE?�|�i�Ԍ}��5
ٌ�74�urAA%\ڨ������{���ld	��Ĩn?�b`�򗋱���|��������k6!2<L��<J��XR�ۤ��cӎ}���N�h���<�.j�AR�Y@��:��0�����/�2<y�8�eYrQ���_r���d2�����EK��R[aC�;�&�r7�ڔ���I�%��nq�S@��F
D�e��g�#Q%�j�� �Z����G��i�%6��)>>��7+�%ϋ���z�,�X���A�]qyt��R̘��v������n1]pu�nh�;�P�h��;�e���|��^��O��$m�f^�|᳅ؾ7A�Ll�L�j�� d¸!�������%�3DI���^�fR�N��������eر����:9_\^'�:�K�f�g]{����F��TT��gO�]۶�z�+3�G�H��j&W8	W����]�ĝ�I����F�Jj��4�T97^}%@g�lzq��d��� '��	I� ��	��{wǢ����L۸Ǝ��R�Vz$����1J�/e�l�;W��_xB]��)c��T3��yIf|RnB��Z�6��_`��,K��t��Q�����Ć��0ȝU��S��}�W?��D�*<-���V:����~�r=ZRJo?�vg��*��n�c(A�r �����n�7����smZ�Q��,S��5�V��ȭ4��t���V��$���P��������Tv�9�|�LOH��(�)��(�P���A�+�7�]Vyf��M����{��6��`/�ސ�yI�)�$���!�@����.�?]siJ�,��T�I)�C��i�aq�	�n|�h)�fLS��g��#�S�ug��^�d�2�}�:U-=�Z�`�ߦ2�"���o\�ڟ(��!����'�u&W}'��:�kM�-9�8(��=l����"��@X��+�ڄ�V��ȼ$�N��D�֣[g���Sٕ�r_�5qb}A�C�zZ�����x��=�����g����x�QU�< �;D�;e󭯜�Lj�"����gaL�89��8�F9�+�e� �
�Pr�!p��`��z̆��lݦ2�;ї�c g��/6ɏ���R��c�y�*�Qp�!��Y��Z�B`�7Qw>��
�Ibs�4��ek+&�\�$�^n�qb۵US*����;@�n���>[�#�_���cY��Ȅ1xq�oGT��١�1��t2r]Fu�M�E�3�� >d޸�}��#�(�����]2i�@�8�5W��ŝ#����`r�d��x:�b�����/��[�߮ 1�3>��Ҏ�0V�'Y��Y�����@��P6�Is-5�L@�_=��:���&[J��Dn�b��@ �,Yڣ�Dƈ���j�����ӓx��;a��Z~+��a�� δ&�W��F�|��>��v�P2ZӐ� ��vѲi��q%60����:5O3��g�g{&�^��ulO�E^�`�{�n���p��W�>�?�	%jk���jɤ+m�=c�1����iq�%o||�q���W~�n�����b�GYR�����?Q�w'��N�Բ��xq���J��xzΗ�{�0���|6_�e���:n`�؛�&�A�L��٨�a��QBw���)y�38L�j��Xcߑ�����k���o�	ǋ��Dؙ4�p`G�_w��b��T�/�_��R�u?�w����HQ�����^���.ao�N�|��E��MTGd�z���.O\/��͡�V��C�_�7�!�}	a���)_��Vn�^����|n�)J ��d�xwҡJK1��=���v�*��������)�ɻ_o�O}�~zK�{�Jb!�M�j���a$�6��^��;l��r�E�&�>��L��v�YY���e�^���K>������b�S��G�J�����ʭFT��S�~Z��g��񮹄�	�Y���,�h����ބ1��!���>��k��Iz�r�X��7�s�s����8#cFeJ��e�\��I��E��l�*p�gNu ��Y��x	ۧ�d��A�5� q@��4/�I��9(-QI7
����-&�P��,g���5?[V�Ǝ^��U�մ�j�7iEE�� ��mc�Tu���8�(-D��bC4�����H��?� �u2�#R�1�MoDZN+l?_�\�u�}�ք͉}���v�i���W� �g�aSR2A��;����J�aOj7�j��&�qU��Neb����CAI#�܏��ǜ��PF{�=��0����n�?4O�&��8$�@��2 5$�Dd�k�����*���M��51 j'=(� � ��PV$e���P����� �]�����xge�zF& ���q�t֓v�v����) ��ad�����Ɯ��u:��s��s�+�r1���Y�m��^A`.����>�)pj��w]GW������6!�U?o��k{��Gk��O!��f2�Gf�8��8���9=���0���&B���an?�u"�I��*���w1��l��FېU��}X��V���Aܱ���2�E6��#�e0K,.�;rG�8n&�q��|�#��	<��j4h58�$��!M7K}R���t��/ NI��뜶��8#�u:�7Uj����:�U��yP6��DԮ��J&����p�)�р���N[M��;\#��2�� q}�%5��bL^z�'�ƨg�ڻr鴆�̎���	�ر?��U��/v&Q�@dy.Etvj�koRn0dp8CE0��?,�DDW���    IEND�B`�PK   `��XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   d��X�Lq�	  lH     jsons/user_defined.json�Zko�V�+��K��%���o���M� N�Ap�	Q�T)*i��ߡ$'���z�.�!�)���{����y�i�'��:VoCLy�|1��u^��pF��z�[���v�ǥ�m�=��&/����+���:�+�Op��y�җE]��e��o[C�{;'�.�q1��뜲��)!0R{d1uH;W�P��/~�ǵ��U�s�������Ac�� �AZ���2zN��*[���k�n'�Cu�)J�a�E*�'�͋��y�^-�r�n|5��[�\Y~�^'�w��)�_6�Qq��*s����:o�/�
a/n~�ק�_V�����6�5K�bs�����ߟ�_tÒ6,��o������腥mX1
�e\Ǻ��a�(X���^T�FU�PE?�hc�Q�?^��l��?�Z����k}��JG���^L���a�cL��mZ�q�J�Aۤ�������)E���)�m���S���1xA�A��g����#a�O�a;8E���%@Ҧ��p��J��"l�9�6��O�Q��X�~�Ҏ�%�����Q��HXӏ�Q��HTݏ���6k�AU��m�Q2U���)�-cP���[l$jB����D��(]b$j?�XG�#Q���:���
�z�mc_��Ǽ�f�wx
Z�]��%�\3��q�rL;��]���X�7ث�\Ū���a�7�;G���i��U����lx�ep��z��/?^g���Ǎ���׹[��ת��f�ﶁn��Ϣ-6��zS�0�gz'��4졇G�"�͝�"����]|V�Nډ�%|]��ֿ���|(�~9U͞�q9��ź�i��b����QJsG0!�e."C$�!�U�k�c����+E<�2�WB#Mq@�*㙤�+zw�JeZ1I�.�:�g������ҙ�T-(S,�r[����ŏG+v�q�}vv�����o��n�>�ޛ���{�xB����FZS��iĲ�:��?�'�����nE�զ>�.@[�b@FX�t-�^��B�����K�G�#	qP�H�Q��$筥·C�`�k[�/`����Lbf�3�Exxζ��Dg��m��Rpd6��x��oT�!O��4r�+tt-b�IPȝ�_�6{B�c���`��8ZG
�i~�6U���]a�<>?I���PŵI�Bx�x�-d�D|b�@����J��{[Pc^F8��7�fF�鷏����������\:p�$���#"G>qƹÎ�������@�@/����q"�I���eLR��+BYi�1�+��H����董:�2�1�bD&9�-�<���	�J阩�g��J0~��`���5��YP��&#\Ks�EW�&:����Ԙ��@�V񰉁UtL��ɠ��f!���2�ZD�TB�L`!�B3���<�	�f8�JbgAaA�l���6�
h�3F��(��F��M.:_lBIƸފ����e��a�,p��g�rh�GM�����8����Q��5r1B�s:0��R���۩�������軮/�k���~�~Tp��_�zV�٫��G�A���\��!�E�s����H�^0���[��t�4!k��	����^3�;xۊL�qn8���hFߍV���\7�X��`��]��x�_��?~Ĩ�C����X���~�v�%��b,<���W��7���טx9`��~�cM��U���X��ׯ���!%O9�H[�D!GJ`�|�O�K���;[C��ԧ�zӆ
.R��X0d��H)u�)� 6*�F���V�K{l��;����R�dp��E�˺�so9�l� �hn�sX!O��2	G��k�(#�t�I���y"aTC�@�[@�p�ᇄ:F�݃7��迎
Ƒ��ߪ�OQ�W����M1�.�%��|�x�=��ޛ6�0����H�9c<J�z���@6�c)�0 ���b����Q6 ���&(�3;�2�<n�HO�A�b!�y�I#���<$i�l��k���sh~q\y�z��Q����n���'J�$���i0$�hT?et�K��ř���l��R�����0����y�.7<�� gh
H����zkn2����]>]� ����\��]�/C��M%wY���ը�$Y˙�����hj�Ũ��=��D��$y�T
����6)����Vy�i�|���eC�����3W�:�&��B~���gu9�!��}p��A�ٿφ�]�[j<���yZ櫳����)�߿��ۇ��Ŵ���wU�)Ԁ�~P���gܚ� �V�?X9���W��D�ʢ����9���#g���jv?9���I�(&�it��Ҝ
��r�'>O|��<�y������'>O|��<�y������'>O|��<�y������'>�W�����PK
   d��X�kƏ�  ��                   cirkitFile.jsonPK
   `��XWC��)�  � /               images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   `��X����7  �  /             ��  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   `��X���a� �] /             �  images/43b8fa2f-aa16-4fa0-a6a4-ecf006c83c4c.pngPK
   `��X��НR5 �� /              images/52cc771c-8bcb-4758-820d-da79c3626c72.pngPK
   `��X8�Z��(  �(  /             a� images/52e5cf08-beef-4b5f-967f-8676d3f3880a.pngPK
   `��XT��"  T$  /             �� images/53cc934f-9b11-4097-8823-694d19808ece.pngPK
   `��X����+  J  /             � images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   `��X��_8
  3
  /             v/ images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   `��X�?HU!  B#  /             �9 images/585092fd-6de4-462f-8499-92296fb2c536.pngPK
   `��X�&�}[  y`  /             �[ images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   `��X$7h�!  �!  /             g� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   `��XXs�銙 � /             �� images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngPK
   `��X�Y`�1u � /             �s	 images/d9bcf815-618f-4ab0-b416-9f611d86ef67.pngPK
   `��X~��a� ٮ /             �� images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   `��X���  �  /             �� images/dffc241e-8a0d-4217-bd54-7504444465dd.pngPK
   `��XP��/�  ǽ  /             �� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   d��X�Lq�	  lH               Jn jsons/user_defined.jsonPK      R  x   