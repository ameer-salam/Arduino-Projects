PK   �v�XiJʥ�  m�     cirkitFile.json�]��۶��W��/�X˗��N�h�f�M������$*G[�:W��t���;�䧬cZ�$؃>l�3�4�83|H�0��[���e��ou�*��䚆�ɝ��wj�*�N��.�+u7��`������O*����y$�I�}���(�~���4a�<�Ԝ������x���)V�3Ѐ��&�;8l?-�ܗK���)�$ɲ�ב����ey���4TTDZ�)�u2���j � ����C4�2hXd.��̈H6��P9�#�hf9�ct�a5�O��
@� ��cexX����* �ͣU 
��G� xW�Sq��9b�&8�cR_(~��Ń'�eLb?�T��ȹ+�T��űNXn��d�A�g1��υ
�@&ԏ%�~��$MT�Z���OB��A1?����<&,�LSf2]���;wbPtj>���8�P<��K�6�5 }C/�]*���(s��q|�T��)�}��-�u${A��0�p�V�����B���C�C�8�q9�r�1�cC�F���Q]c�F��#��3V�����3�`�p�VǬ1Ę�9��!�j�����Lbȇ�X~\��R������X��i)Bs��P=�3+�a���H��h�$~���WY��Q �J�:Nh�J|�u��6ܺe@��m(�Z5=��Z��>�w�jyx�XN�>�8��q!Z��?�+�L�0���q�'������	N�"����y�֠E��D�5��n5�����B�HQ����#E���D�5�}n9R����A�HQ��Q�(��h�!�]!r���os�"�ymwnۙߦ��+M�Μ#L�|7u�]ijw�ar濩3>���=Z����{�p��ݾSy��;h�����z�.�-qlĞ�5n�;��GlD�P3�FGlK�P����i�dpS7,f�t�9bi�֠f`��zC��&�84nX�ܰ��a1s�b�Ŭaq`yӰ�汢&�����/�ݥq���s�/��v��ζ�q`����v�Á��|���p��,��Z�F��X��qd�E� �Y���:8�rֿ��l�naU�Z;X�_�u]�~a߁�va�	"G�څ}'�)j�� r��]�w�ȑ�va�	"G�څ}'�)j�� r��]�w�ȑ�va�	"G���}7.ҝ�v綝�m��q���-����wSg�ە�na�&g��:s�C�F,�����x-�����2���x-�u��>^�@���@��9�1�Ը!�����@�S7$�nX�ܰ�9��nX�ܰ��a1s�b�����37,�nX�ϲ�za�����za���p�^�P���>^��>�^��k9��za����ܵ^��k9�]���X/�㵜�#�����S���n��ϋ��䚒��]Q���~�R�͋弬2]M�_b�CE�WS�#����iz��֏r8M���3�g�Q�6���-ؿ���k����l�sK��Q����-�
&�`Zƾ���=[���x&bZf����_��W��Z�7�[�j����/���L�(�h�G��x �ػ���ES ' ���.�0.��%=x���� ���'��m΀�L� �aܴ�y�j���i���m ���u���~/�|�=-�.2g��S�(��@$
���L 9�8P'48�o)���d ZE{���=�D�Vў�C�@�hO��A'4�8�1�Rh�y?��s�y]�^��9��Ł�ѝ���p�a���ѝ���p�e�7��1�lF�7NF�����x9�ޑ3�$�a_fuK�	>#��a�!�{Af�a<�,]��x��;���s�� �s(���D
5�Na���ș�n�A�#}{��Hj��b�e1ò�aY̰,f'X�Z���P�c�-��Z��ȟE������}����u���;���S�wp���[���?о�;��}�>e��s��C����=Y�����l;����wG�"so�����9�_��s�l��k���8���I�L�bn�p�d���T45��JM]j*SS����ԧF�	f$X��H0#��3�H0#��3�H���6�j>(��/; `�l8� D�~?T`ޔ�n�y�k����Eٽ���=��~@C�0�f"~��f`r�9�b��[=?�zA:&���{����?�<rڟ�a�y
�����>?�;0�ϝP�k�<��߸����w��6��*�O��d�Tמ	A}���~�X��wE�_tEA�(��~��D�HvE�_uEM
�����e^�Ū6�c7j!��?V������x�/�G�|}o�Y�ra���M��tS�����d�o���<`�U]��`��zc�����Z�ͷ�Ͼ�)��1�zY �	|Zݕ�-���unPA�JW��"Y��J�k]T:�\��Z��ߨ�:Wi��t���j;,/�U������n�rU�ͯҿ�E!�	�,:e��(�bc�( ��O@�$�S� ���f����Jk�	AdDT�7kk���]W��%:�@�^�e�*�J���*@�j�N��AwQ��u�K�Y8e���n>G$��"E�����z�������0��觟���߀F�W���v��ȧ��"NX�5�4 ��L�[ǹϣ>��S澦>	�u�9��R����yY�w,x�3"g�>9�)e!Pǧ�Q�lJ>s�f���s(勉Ϙ<��S��4�kp��i���C���ZJ+�XMxG1FNa*�aL�|C�C�(�	*6Y�ԏ���0�h�Yx�K~9�}"���4�>�֌���NVKv��c����a�2e1%2�P�;!6wŏ*D���$���]�x�j�8���È����|p*�ƶ�35ڈ���}�Co��E��M��D3I�x�ߋ
��T��&��a. 2�a�T$y��yJ�^�Z��b;k��1�0<f��a;V
1#�ш��<��K7)0S����f�MMiƑ��^�=]������5 �G��A��[[���<<��N�������Eמ(v��f�������k�]Ƴ$�^�%E_,a�%��P���Z�wi���)ohl���F$��$�#��ui�S�9��Ϝ�}�:<ػ.��˽���:eQ�Qb�+v�BK}�R_d��;}0���qK}��>���O��z�������
��İ������vf<N(�4/���n�t;������uzw;��N���ъ��3?S�	IE$�B4K�4А]4����E	n����I+�b�a"��9�����q���qB�Ԅ$��iO.��S�ܗ<a~����(��L5M��f[�'��u��(I������T�WBG�Li�DgQ��\=Y>�F�/`�ۍG��ɣ�b��JdN��0�~�2�4�e*ɹQ��@UUY?���=-q�"-i�`��(���a&��s���hQ��>H�H"�G<�� 5$:��$�2U1�ģ���߫e���	p�{��{����_ɲ�\{�Z����˲ޯ�tÒ.\y�=}�_馬�ﲬҫUS�b4����ӼX�D�]3�8Wi �C�����lqH?����xvd�={h- �3!F���
��*���9qΡ��Sd���3$	�-��9�� �� � ��_H�����&9iN�C>L���z;��X��u���zQ��;U��*�bv�����^��ޖ�E�'-!�zŲ���9�y����c�x�����\.uZ{?=�z���ե���b��_7�����0o?�%���eYߵ߯ZD�N�׍����x�yf����Mw�ܡ��e�|jA�Z{�[5�e�?������]}���(��HA�ؖ�Ò\-�rXд����e���z}���.x^�I�~],�bH����z�R���6��޳�~���W�D����)�L+�n
��{rF�WY`s["���%�������{���[3�T]���js�Y��)��;ݙ�nio����5>�YoQ�;����cq�VsW_ojP����4z�F-��]׺2�!=}�t�䕝xz�*/��<n��嬨i�u�by�nv,���[/m/��Ƚ�]��B/_�wp������t��o9T�}��w{{;i��;��촁E��E�TE�O�����O[��V���t+F����4j7�?z���@����������H�-���e3�Λe7��bu�e��3��Y���@��Yf�*����i �1��YKl \d�ټ�����{���I�TL��8�F�j��b��u����@�`�ʛ/1T�Xj��s8;�M&x
�e0���ŏ?\ �xܱc�fXPc�"?.W�3�Yc��!|���E���O��F0�v��!��^0u�v��S�	C�U	�Wpa%�H�&�/�r�m6�qJ�,
�)�S��{�d����@���U������m�\��9�$����sm&qb�̯TE(�<� G���呟�f�9��M
B�˄���9�9	S)|N �"����
@P���@X&�}�5U��&��gs$��x�kJ����E��]��Y��X��P�0�Ea��^�B�usM���0���3����ݵ;mƃ�n��V����߇��	IH�t��v�����������b%���X���;�?��XhU������ky���ew<�QU�w/�b�?��w_��Q�]��C���g��)h���\�~i�۬�l�U�<��!1����Av��[�^}��4��۟�s�瑻>��<r��|T�����}~X�pok��{�N�y�Sg.�<p���q�N{���q�5��㌜���Z��ZA8����� ����|��.���� ��.@w!��vH�{���y\�g�{ݿnWi�fv�=K$�;�EHv�/J2qrXp�B���%�ӕ;r�� :r�� �
r��	rG��I�|D�Ã;{1n��ωZ�c��;�s}.���������P�;�FO��?�%���fGڳ`t��t�;����v���:��5L�����R/:�8�N�D��N�7s���J�	�i���ى���������$<��G֋]?�D ��$�Q��΂F�ֱ�IW�'�A2�ѸO� �[&<͔�qK|�����Z�\�������ڵW��0r
GՂ�,h΄^Z�̈�5��<�R�xB-Nf�pu߮�P
*�Բ��֐��.gD�c���`s�p�Z7>z�bxNtTm�kp~0]��e�t�y.ݺ�3v���؜qcTZq�\��s��u��E��$�f[�X,�忨�9T��\:������/j�V���7Oj�Ɯ~������PK   �v�X��(��8  �8  /   images/02932828-f6d4-4923-89fb-67d65ebd103a.png�8!ǉPNG

   IHDR   d   �   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  8kIDATx���T����������tX�,�(HS�(c��5�ؒ�1&�3��&�F�1�?1Ѩ�1��i"(�.,�l�;���o�웶�]��|ٙw�}�s���<ߘ1cZ����&�x<��z���K\\�466JKK��=!!a��f���f�w||��{���!x�#��1��|>�< �\�r���>�v�q���͛eӦM2e����dܸq2l�0ٹs�����	��}�G�ĉ���J^y�)//��=�IIIr��'˜9s$%%E;�0ٺu��q��.�E�u�(<�]p�:,��g��:9##C$999�x�m۶Iqq���Yd��=z�̜9S���Z�߿����K����g��C9������'//���'�0s:T�-[�_�y��Jee�A<�~��f��ٳG.��2Y�~�����KlϧO�>2`� IKK3g�޽��555!�A��Ғ��w�O��Ө(P�6rݺu�t�Ґ���v��an�U�J�ٳ�lٲEv��%EEEf�u���Y����3�\\��� ���s�]�}�v�����3c�p�n�4i�2��Z���^�>r���J��/6���gAX��t�0ax�R�%J9�t�$(u���Pޚ�������_���:�\��B���w������a�\���ZxFvʆ��n6���q};Vw�%��W�^�JAAAȯ���S|���c�����#	z��!cǎ���z����iJ�=�!v�#F�xAW��M�� 7ʶ}�����o�'�|R=�P����
�%tvn1+Y������� �畕+W�"L�n�,�e���V�Q�������ؕ�;,11�E�[��r��p)�*�B	��-�N�����P�W���9~�m��N�ͼ�_�כ<���
-���?�8O���h��TU�.��w�q�lۺM�9��y�	RUY%wnO�
As��>عc��=�9����o��V`��+������J�,^ I	>y��G���e��r�7N�Q#�ˋ�?+�e%���$��		�fa(^���_���%�w����7r�5ט�7��>K�K6� H�6;D���}W^ye��gϖ;���S]q��΀Ҭʐ��������<�w���eM��*�q���Q�Ƀ�Յ���&3$>c��dű�;�H�lʢ��d᧋͹��\I���y���/iƙ��v�_�w�<5w����J��������7�IrS��Iz��́����n��{ｆ((ʶv*�W�=�c��y<�ET�3�^8X�A�W�ҴZ���:�h��47���5�����|��/���S��رn�(���o-N�#�:TD{P$��߷�rK���.�j�>S[[kvKT>j�js�bn��|<����5��Zb�(��s�D��Ǽb�]�yc�ӑyU����<+,�9cΫ�dT��?Z]ǹ�����;�4�n��V��+**233�#��i���|�8��$:�#���A %H��<T� ���Ȋ��KmE������"i�x%��@��;\�S�Ϯ�x�i�\�y� q���)��=���|�^�'i=�IF�A�OT6�����2���U��%ez��U��KL���C$C?]��MQ�G�EM��Ç������޽{�sss�a���)!��Y�Ǒ����=?p��G�e���u�1%T��Q5���]��SZ�S|2�~)���J�����LK���ee]��|��t7T
 �-�d�s7If�Qr�ٿG���mPB�{�ϲo���'�Jz��뽪*��I*<$���Ȁ����؅�����d�+wI��)2�?��l�����3Y������Œ���z�U5��a^�T��e��ߓ���"m[D��[�r�jY�R�}II�T�6��a]��t���O>	�!2����������<�4��q*�.S{dȼy��;J�/QJ������L헱��K��s�qSJFZ���`�������u�����oB�C]���RQ�.�L+�Aj���ŏ^#Ǐ��+�"#�$9)^�A�U�2��5r�_~*{t�#ξI�g�aW�W�H�����#��Z��m�+����3��"��d�jƏ�"%����ܵr��W�ލɘS�	��V����by���� /��1N�����0���s�ƍ1-��7L�q�5*;??�:%�uF�c�~���F�t�l�ʽ[d�?����)�~�̙�A��_��dמ*��'��8Z�N*W^��,zl�L��{%�N7kX�]@�ؚ�BY��������՗�nvqCc�46���3H#?�l�����e��"�}kP��Ƹ�V�;NO�d�+��;gȌ�#���IWs�ޯ�k�3S���'ɱS�ɅW>*k�H�Cg^e�+7��P9�}5V�}�,|d><�-�!!  
��+d͚5F�[�X�s�GV�p�\|Z/��w�HUu��`���x|�Kj�z��F����˟�8KN��aټ�e_g-��Y�>W�x��?#U���t����X��#�u�����o�>C�\����͑�+���#�}N�+e�[䞟-'��_��o��]R]� �����>SN��)5Mr�n�� W�����Ø
(F(EVku+FQ%2�V�u�r���l�XR*��U��g���푕,�Jk�fq��J�F��x����صߛ"���w�a���(ݱN�K>Tb|��Pb����݉�e��WL��zD���}^e�;�͑��r��ce��RIJ�Ib�W���o���
��/c
�ȅ����T&_pgTcֺoX�����m�H�ٴy�"����2u\OeK�RS�h��#E�o.uv���2E\��x�����c&��?,������
"�UVP��C9�l雗��v�Ab,ئ�n0��:i�yґ����[~��RY�M���z�{?}O������ҝ�7r#A�aR������Fe��N%��H��
�%�>?�(�����!��&+9';IW\�Aۿx_���K���{fF���U[H���2�G��f)��kŋA~Y�Ab4b;i�A ��/WeZ�N�8:b��F���)���Fz�<��&��Z�+��jw��8�i^��=UR_]*��i��ϙ ����M ��� i�	RV^�ȑ}5F{q�0��y؆�����o�x���vC�r�Ttb����j�So�[O�Yţ�L"R�qd�e���wX��7G�����;�c�9
�)��l�X��I��'����d�`w�d%Ii�#GXٰ��D'�V]S/{�5J^f�!�X���Ȗ�k���#���Ęf���� nϾ��̍�@�y�{J�^�r��CU��5;ο�@�����/��+�T�iI�Ĕ���q�All!�66�	՞�gw�1I>x�ߊ�:=��	#G6nq��p��~=�)�͖��G��[�ad�{�)QJ���I ��d�V�]�!���n�2/ZV������K/�dvq��18��6�\� �3D�y��ﭒг@R�bz�;
����	a�92HTb,̶vJ��Qr󏐵��ǞY&W\|LP�쑝���k8���T�?�}�����'�EU{q`�6N>xs������q�!�8v�@e��Ab����:o�ߒ�䌨;�Y-�AGΔyy@ޝ�Q��rQ[�<Σ�q!�3���(�W-��!3���"Db�˗/7n�~���D���G��)SU��N���~�%2lH��x�H��X}i��F+���*O@�Ϳ{M���i��g�Dod�^ϼ�N�_y��K%;;U���V�-I�NB�x#7�r۽o��M�2튋̼�1��<4���W����z�����a����Ӣ��IP���R��$�3j�s�q�ع�M��(";��w�5���1��s&ʇ�+T�M�|�=�6�䆟ɏ��K.��x饚;���o�+�z|���6K&�^�lV�k�1o�ae�)�����1�R~z�q�B���ei��?�#/,�Ȥ���80ٹ� kښ�"9���W�LQ��@������a���r������t�/��q0�]��u�WO��ɓMX�
�j����c�k�-�!~��������-?��L84K�A��(��={kdgY�d�<U�~�ʪ҃H3<<�^�g��e�A�O7���]��'d☞2����k���5����5����Hbz�Qm-X~�
�_���~ ;�����O�}p�Y�#�z�� o�U�e���s��e��s���B��!����6�*�.���a y���c.�����TVmZ!�%�ū�+}�9jȑ���� ݽ��i$e����Kzn~б螷��{����-�d�ƥ�֢�FcJ�/��3ɸ��m��H� �9Vr��s6�K�C����Stޕ�p�j�_W">�aه��)�����&\p���I��w�.��]Ch���hH��5o��o��0ZZu�f��p�sN�d�%�.��1��*蝘�Gz���~BH�ə72rɽ�:QrG��6GecD<�1gވ��y�b�~��!8q���®`G����x���!?D�TĘת�!;"rq�o�і� �yc�3os(��ɶ�����,Q�z<z=o������jYhP�����/���Ӎ�E�	~~��a)R�v���E����(q���^��� �|w`�d6R'h�[�*B�6�9������!>���3���o���  y֬Y&I�"DCT_~?��3C��_~�e�k|q-��{���>������<���Ki�A�cSe���ciA�x�bg��xꩧ��N$�p�Q��裏9�q�Fy�wė é�hb��8
C��;��c���ůApjR���7K�����p��/�ɲ���D;�7E�Q����^��J|j�7�oSF��!}����/�-/�چ��d�z%��(M���)��֔G8;էc=��c�H}S�|��"b��_r��Y�I	q��Ty|~��'5(�N>"KR������A���2���*�|��s{��Kf�7��U�9���	y\����Izr�؊Z���b|��+���D<u|�Y��,,1�fGI���N��u;k�9A�"�oR|����OvD�����+.�
�A���� ���Y�Z!ߜ��hۊ��Uef�����Se���^�j`�D�')�����^6�3��=vH�D��mv��\T/[����2@L�Щ���;����ʥN�N��}�y�N��t���Qį�V#��$^��6��������17��=L���k+�̱p��),k�:�����|y��r���ʱ�3ewY�4�[��D�����d����g�HB��7.5|�-Z-�,t2�T-���|;fJ��i�qf�r:�Z�1��}�RX��K@liu���b䎹%R]��w�V P ���c!pM��KG�׉���qeO�yڮ7d��-�+�T:�_���JaSd��dx^�<��^5�[�`��v��� �����)HX��u;k���c9A��� ����<�v,�\e��x���;K䝏ˍV��/'�9�^�Wf�a[EM�k_���%�D�n�wV���"�Kuek�(c�`��݂��sXЁ���,�3�$O�VR٨�ϰ"V��χ�~����nWM�N��0&S��y�҈�rK���ݶeo��M���f�F�o�,��Ň���O4i�6ށ7��؃0�X �6,-
�@�HeQ�Zv�a"��.�!�Peez$H�Z�ŕM��R)�j�0 ;��:/,n��}q�>٧c㾌;_u��=�g0ySii2x�`ٽk�,��m�)�ѠN5��gL�8o�*�^_Q�\H��=��A��פ��}a�HGE.���ms��	b�ymy�!x[c�X춋��Dbˬ}�D�����t��ҩ ??_vn�&K� �A�u��1��'�Hz�7��dm�]'��WF�q���c᰽c�
 E�,t�
b�]�z�!�������-Y�dI����s�1��t<QE���铝 /-��� PO�'G������w�����~wbY�<�B��p��4�����	��������5t�Eň#�����)�h4��?hA��x���Z�I���Q���F�N����ފ�#GP�H��[��t��T*�\x�&�Ǉ�E���_��C�Ô��q��E���)=Ϳ�T~���)Ƶ�9 �;i��4)S�m�����~���:*C��
� ���Ͱ+`Q�k�_z�%�e!�����,N��ɥ�^z�����T?��F����k+Je�jZ�(˸ٱ�Z� ���6��țE�dD�d�^�a,��D˲�������׾&�<�1;(4� �Un �$\�_ a�wךh��w�E슺�f��o6!QU��d�aCᮓ�6W��?�Q#���F�ފƮ���$�m�ԩ&Q���g�}V^{�5C�0�C�������8bH�	}���Mmz����V�I��ũI>��iʆ>X[a��l6Ao5 14�-J/��U[��;�m��� �J�޽{��ˍ>����4�>EV{�]���o\'9i�&"�Ya����A�a��_W;y��FTq°tc��7u���� {�Du����!�	'�`�`v�]�$p�� <���{�VY�&h�oeC�BeƤ�Fi@y���ii�.��B Mz �%�<�Z�*�P_A��A�����e��bΕ�P���������p0Z/o�ʛ[��<��kd���6Y9�,�E� w��/� 6 ��&���o��8Ot�kdA�,�Tm*sd��4)��aCh^�J5�c;'�Xe�ʭ5]j��b$U�Р��H
.{�A�zx��ϝ �bx^rH�Y�\�E��l��=tGʝ�4�U6D���I_௯,�)�g��66ICWʐ@�������3�qKM��?�|���,+V�~G�xx�	D��xB��q�/�P)o�Ժ�]��į�@Ö�u2�"��+��x;�z�+wrb�a���W\a�	���'��~��"�����J ka�s�8n���W��eJ�W��H�����yb?V�w��&��������#yJ�:��r�9Bl�8�!h�C�&|�nۮ��pH��SO=%4�a�!*A@.>({�UWy\�=�9�m1(��x+�A-�uҨ���+6ε�a/GI3�E8��8ix��O6A�-E��dO�!R4�C�����VXTѵZ��#���$^d	�N�������V�ߜ�D3f�0:5�0J�8�7��_C$W>/����T�;4Sm�����Ę�qy��p�z�if�%H�� d�'7���:�Ⱦ�f��ۘ�߻:/�P]�~�_�n|Ʊ.�&x��G���r�6Y`�jS����G�L�/5����$&����� KA��1z�"-Z�
G��;��T%J/բrt�3_a�"sW����~9�2�_����u4v����+��X�:;�o߾f�����i��v�te��5��v��`V�*\�XIZ�Wv�8�`&K��Dg<�jXRhB?4U�	�l��7���j��
l/i0�t蛪��jv��Bm���׿6��/���}�٦0�̰�o��4}��H9bB]���#z��o��b�X�P� b[F���S�e��Ϫ�C)D�<�'K�&��OV{�n�z��ޙ	����bR�
.uv��nM��I�g��|C��j�W���Թج���׿�e���v�i��B���QG%O?�t�	`���`U�$�b4͇��Ak�l��3X��d��&_������l�ߐr��#6E�Ly�G6=�N���~]�]�Kl�&�Yw��	P��!�C5��&b2ā�ݸ���y.���Ξ���,Аȟ��C,��!ҕ�Z�Y��C|n�CM��RGf��6� 	v�8���Ů�,rT[3Z���O����t�R�ԅ%�ǧB�v�DC 8qb����:a��r���,-�=�fţ1���0��`m�0��cL��d��GC(�� ��"�q���թ@�8G�?���r�uי������T/êº:�C��
���O7�%���af{���`2d @T�'�1dՃ�}��mU����O�el7ۢ�g��tY��p[���SM���|`ކ�]bm�zWc��b��`:��7�鮩�
���������m>.+�,D��hP�T��)kPA�J��v���#�EL�ú�dk�ݠ���[���v�,��+�m�(+((0JS�XY��ّ������{g���a'~Za�%���U[�=���j#kI�ț��V�1��p�WWB�l�r�{�����$�6�j����Im�u�=XS��E�z�hCMK�aSM��C��@�	lu׉���k��ӛ����x=��=jQ7 ��x:�[w�6_yp(Z1��	p4v�mj6�W�.��'O7V�b�I|q_"�'�����&>`,�i�B���iӦ���~!KȘ�-f����9�,�]���h���� ���y�xĿE˒�������w<넁8��w		t��w6��-�Ƹl�m-+���&����T�v,��]��] -�^cx��e����i4�g�ظ0��}&?����,�lMp�E�����F�W>�L�vZ��΅��.M�ˌ�n�y���Hqe��+�ND��c�>����}Yx<��ᮤP�`����m�56BC�dkjM]`�4L���� ;X�''���J\�<�JEVzs��ek�]���B���D7�K!$���3�L�O"�c��H�ƽ�lm'#q��d�*��,ͱ�!�7,����	�9pRw�pX<oر�.�}�!dH@&�w���z<�|�ȅwה�5Y�!������RS��a���\��0�.�<ei����.�/9o��K�/�$�{�P���4&x�ǂV:�!G�H{Ƣq��.!��{m�_�I!� i�x{�����n��p��`�I�t������ԟ�����$�ט�	�o��¿��`ߤ�m�����E�Ŝn$�PI�h�Ð���%)�qR�
PA(\�+�և8'�H0;���$�C�~xW!���2d.B��¶b�V !|�&E��>�������� ��XI�����C�����o����>:S�\P,q.����lA�Ӄ7��X�ZSx,�R�w�{�9I��V�Ww�#�����BXԨ�,z
v�$��w�$������]l�F1l��-D��LS�X�Dd�2'V���Ǫ�k��;k����'c��I<c�;������~�9D���5�6w��Pv &y衇̿�Xz4���<�yYT6��Wl�1�8�:t�|[92� C�ߴ�0v��Ϧ�'Ȋ���M.�g���Tn:�B��?&~ī��P/��îx����N�,`[!�݀��7��w)E����1�4P�+?2E`{q��V�k:9d�U�_[Q�dǻ�b��|-�f$�� �S�F>�Ġ����f��զdAc�˟e�� mX^��d�����.&��O����|o�Q�ρƌ-S���QwESk��n�#C'���Z2≭�0B�o� �$����k�4��x��w�I�c�G��`�;���R��-m��Ml�D��_�u���pv��:+�DY��
���"���h��:��v����������� ��u[�P��@nG�u%X�XW;�ŉ��x��fnl=_[t�=�6���l�. ��8a���Z�C�䴁g<�wSM���l#zsP΋��`�0L@*�M"�z��
2
Wms�O|����A�;���
r�P� �]���%���	V;�(^V�0L[�X���ɟ��'�$G˾�
����o6�YQ���j]�:����,蟓h�������^|e�-�}g��dD_��Ѝ�������JJ�z�}YV��\d�8��sx.��7��Ұ����~����\�gN�a�uV�W�\]n¸Ѻ_��N�|����f{M���;&��,V?�E����vc!���j7Q�=�����o�&y�^(AL��D�)�yn��R�~��=eцJY��ڴw�uB�W��Ū�� �WB㯊�%`��*~9���i��<�m�s��`S�_~�! �qd,��?��pm)V8ķ�e�9O����������:"K�_W�+��$���J0)A�+�X	QB�`�B�:*9���f�,��)��b�R����#�Mׇ�n�[��|�?��O�;��E(�`q������t�����R��g���cOd�����،Z���C6�ݽ��=TV-W[�*��}��D6;��d/Z-�*?�<0<� ����;T~yzaI���_Hn�(�nvRLA6V=����-���AHV<,���u��֭w5X_�o� ��c�1,ş��e�������'�:�EJY�J:��^��Vk�(M6�G��B�2��S"���� �2L���r8lZ~�.���~� �����w�qH>/� Ų6��|��̙3M�
q���7&?�	7�tSTyb�NrA/,�ՂgFXP�s��qJ����%��#�#�ߑT�����Gf�U�+�7Jr�	(I��%��v���!;�`�P�ЮP����?���L�ܝJ�*Lw���p iu�4bqr�DZ�-`y�[�a�õO8,���+��-��>IF��;�p'Ũ;hXoji0���x��z������`Kz����TиPy	\a�>�q(�/�����ch�A	 ��Z�D;��aD.q�ʭ����h0�!ׅ��?���^{�r���{┅�G40�l#�V�uCa����E@��� ��|�»#E4����
{��z�3�zDT�L���J2(�z���`;`��4�[*r��⻂�c���M��n��CU���8�Bk$����b^��:���z�T��[a� ��L�	�/:Б�� ��K%p��!+��HU�_��2 ��!q�����u�����!��C���i)��w�)�AI��\�3I�q�v���I�&9��h2W
�;݃�CwH�dAr=2��*$X��U`;ʡY��G�>��!������ �d~����"��[Kq���x:�Vo4)�MF�#�Q�I���=g��4+�a\���z
�J��(�tw�sw����fL�PB��G�駟JqQ���^'�a�+�Z��m����~6!��+`��+���o;;�]A(�gzp)���np�Y�29܆; �0)u#���P��kdO�Y��Y��*�b��7A��7�4�����r2����<]3cL���-�����o�����M2�n(sx�����3UgD�#A��X�$~�Z��H�:ݼ�1�0�L���	�$����.uH�)vH��5F���D9�= ٰ)� ���ļ�n1l� ��d3����߲i���47��Vt��c���pD҈�ҍU!Z�7Д̨�^'N�)*k0��`��w֔��v��N���v�!m�	�����闕�0Dj[��rt���;�=���pʑٲdcU�1\ t����-��&Y�&�3_W�+ٚ�E�(ma��6iҤ��B��
� =)@ H�0����n4��`Y�nք���&;�E�����O���Nt�O�"�.�	fB��K�`��IT2���w^0Sc���t��t��-�u��K�J�k�"�	E�g�u�>$<��Nkw֚RU��!Ć@Se�T ��^�:�N���;��|�ȁ4l�R����f�qh�x�E���1/z�V����ɼ4� �V���0�9�͜��e1���6x�(c75���cu��7E��B��9�F�H�!�$<P�jGյ��!���n���������=���Bڏ�3�˻���\[~C�u�RW�}Rp�p0;{�ؘ���i�iJ��h�!��.`�3�kk	��t������ç����������?Op�G�6�ڲ�X8�E;��S�ۉy��sQB;�� ��[�����ilj}��RR�Ȥy�����벮d����Om�\[��VbFgǒ�F��X��JQ��,"�L|�qm!x5�$�KCRRR�^�DO�T����'��r0��Ma���w�3�y��k�KQѮ�;����l3v��n�3����W_-Y�Y��ܹQ�Hj=�~�"��?�P��|�56+;K.��"s?�T�_�|��m������7�a�<l��n��D���Jq�[O����9��2���*[\ �b�)E�DxVO*ՁiJ�F�y[NN�T��Ew&�JZZ�uw-�7��ǻ�yw�;��n������ӷ��y�Y&��M����7jēE2$?_�y�9���/͑x �X[�y�̙m�Yބ��hԿoU�?���[%*�&8����Y`�w�!+����(׭7K,vɐz=�Dmm�|ec�&L��OG��A$�G�p��	�| cC�h�� ����x�� I��v|B|̱�L<)QbE��=

Z����>�r�s����}uʔ)�_}�U�k���)���AN�Ȉ�
�ڮ\�T}� ���Z�J<F�]x���|9!�r@q�/E~�4ü뮻�:]W�lYү_�Dr|6�DiP�<r��1 ��C�@S��J�B�)}��:P��ލ��ڇI7��~o��������L|^c�������<�a��(Q�Z�飼����u>��]��������q���j%H���>��?m�,��񇑛d���J�A,��:.-���uXEQm�@�䣧���i~Z����t��ȓ�L��4�o���L6M4��L=�p
�yْ%R��H��k(!�B zø���j��`���^�'e��z�=d-���%�j9<i.] �c��c��l��p��ז:p�v�9�����c��Y�<(7��"[�6\z��6oR�۲cG�Z�>b����a��ٺO��k
��L"GF�3��5k�.��8����}�ň7|���6x����{�rsH �M��U��'�b �?$d��(��\��O"{���N��'�"��߼�̂bAd�� D��o�86(�����bR�k3H���hK<0	h������f{�M����L����?_����h�����s衇>AT�7I�<�0D��曏�gK�(Rv��:CU����SSS_��� ��I�2o#��DA4��JҘ��~���7�
�A@������a�}�"�.�}B���� =B�O���l�~b�7�t��7��A�%��6���x.�3�-[��3f܊������.**���c��`^;��IЭ��^��:�c�٣ǲ�s����۷oϡg ڃ�E &q1�R�~�l��ްo�D�Õ�g�,�Y�f�����E�O�0��)�'�	�#��Bj/���XA^��:���[шY�j] ��g�x�\�E�\嘚�(q�����ڍ��T�w�����>~�a�����n�՝oP��	�:0U���"���^��ICYE��lKX�;c�>����<^[ K�=���3�!|�q���ܰ.x0Z	�x�qӥo�L�x�֭�`ڥ߻\�u~��{�9�d5����e�`��W]e
1�O�S2��P&M�l�s����:|�OԶI�{O5����ȸ�ɾ��ED���1c��{�>37����S����N,Q�fԇ��6���@�=	�S��֣U,l��`_��
?묳̃�7�Y՚�.�f��#��;��ew.fơM��Z4��-��m�b�y�7�P&Ƽ mlm��a_[�w��X����^����� G��>3�S�e=��S�>m!Da�^�ν�xFp�BR�'!�8»U��X�p�Lȃ�'uoyV%+���ʰ�`�Æh�ikYm�$n��p  �@2Id��؍n���Jq$���������ޛe��ܯ
�q����]�=Hp�柬~[�a�"c1��n$�k�FN� A6���^�wV��31��@�� '�m��9��]�| ��j��f���ժ�zN���w7����hv�U�16>p�B��&��}^o`�/0v�~�u���h8툽��� �u�嚶ȳoR�����[�B�t�uy�1ʧ����Tu��3Ϥ�؏^|�ŧ��8�t�6�f���c���o��\��+���cC
�u���=��L��e:�P�|��7����M��`��f$�8�U��� ���3�x���u�H��={v��D!�x��Ǔ ���ĩ����(!c�{T=�V��y%z���_�W�}г�}W�ࢋ.�")Ĺ�+ڃ&���UbD�E0G���� �`�灻/��_A��A�|E�n_���W�f�A�|E�n_����[�V�Ax    IEND�B`�PK   �v�XR�\"# � /   images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.png�|eXU���B��Hl�"���H��Ҩ("ݢ4H7X` ()ݠ�ԢA�.�\�t�4��Xx��>��o���9<g;Y�9���1Ƙ��/+AJ|����J޽� �9����m{�\�y����-Iţ��zT�5����]5���&�0VT��ԶwTm,lt��1���6�u-��-����`0�0��o*:���l��b���/������q���<?J|��yV]"l�G��ׇ��?�8\���ʹ�>��N��p�+�{�+�=�������_�~����R�sK��0hb$��������!]�\��|1�����q���q�.I?�_�~�L𿯕�pZ��E��G���;f������!
�|���X|��`y�<"����F>�������j��Tv�q���FD�=t�{�\˸U-��k�V�NF+p��G�ڗ�+]�(Ǵ�=���}%��|�tB��I
~9O��K�\Nc�u�������}�������\O�D�[��oԖ�����
����}Hs�ş��r��8�\W�4�DUTT�$�ns�nľjܑ�����{��b�i�:0g?�cձ<V?f_�fr0C�U��q�+Q\�~;
�c�#"]�%�[��6�N5�]���^֥2��e�(�%�w����{:�{0��՟b��X�Jh���v���Tj:"�pn�G�=�`�?h����M5��AÇ�a��.�ka���i�_}����4�*���硗y�%�ڹ�m�e�T���S�99<�cS�0+̼Pre�Q��r�:�:��V��R��\�~�i�`�KE��Zƙ�t�^d�n<����9�﫩�����x��Z��?u���.q�J�<��O�C��~0����1���vk���I�q(Yih)`7ߑ���S��cf���{�/�n����Ɇ;� ŋ�������M[����ϲ��r�Vʨ�4b���9`x�G�>|8bʹ/�8·Vp�����T�]���G�]��VK����rT�:,������m�i�;t�(q^k}K��DZ�os��X#|���c�fL���YF�;�,�rg�DN�d���zz�	�����_t����?6����x���kf����^�r���oTЇ~Vj[^��&2X���������I��2��!JJ~��gW�v���v�3�Jì,���y��%�K�g�&)�����X�R�o��� H���)�@��E�E�8�~��HKZ���*萞�����l49�!��yRN(F-�`�Sfjj��{��=�U��|-?��ϼ���րo�.�m�|�1^��r�4kf������t��7�\�9~��)WY�j�(�l��1�����w����;�q �`�q9�Sz̤/.>~��u�FX@�w�QJ�$>t��7��".˄�ّ:��I���1�m_��.}s�QS[ے�_����.�U%��QO��7��#��.Z�~]�͐�Z��_�^*F�g�;��O2Z����UWDE-��֎���O��|�Jj��2��}[&�ʩ1?T�?�ՠ�E�}�'�\Ŕ�m���5J���4�6�xJJy��]��z���A߾��uPq:'�(��f{�Q����n�������j���&-(���w�{��VJR�YH\��CE'��q�#�%ڲ�>t�;V���4�c<<N~)�bґ�DLJ����Vo�M�̼O�U1͜y7Z�k�f����	��}5�{���t�>Œa1X��h�VQ������h"�`m�/��ā�yb������]���Q���8���V#.�Xz�Y�i�y�~�*�`��f>���B[9�(뇰��{A�M����P���gy\N��&I1���2�~�R�?Rv��.�λ�jZ��C8u����lK�E#�!������3���D��sɁ,*̬�h7����젦u���ʥ� ��?��a�����]�g�N2ʶ�l�����6�fp:�Q�:Uc02���p���j���"��������ǔ�n�|���v����o����s���+׮u/_p�o3�#Ͱ��D{O+�������^���]?�P�Lll��K���z���Z%��3a�	��&��v<�)x�"b�԰�-��*���%Ǭ�*�y&J<�z�6�������qj��sv�B����P^� ff��tB���122�7�A�]��=���t���k�`�3MCIK뉔��]��� 6 �f���KHH�̃�����X�S!�K����]{�UHZ���c�D�b���`��<�mH�0 m�֡b:���U���3�K�$������_�8Ե_��1�@�8D�V5''�ߙ�e
m1n�}�����ҧ�����w�+���9ߙ�xո�0�����ry����l�B}0Gp�T���P�t�~7:�����S�6mfҰ� A��c��������"��&���55S���'�"G�f��M;S�mms���0����Gp' ���g8{Rղ���o5G
�t0����?*�G��_8�fa��W�ڟ���B��`8���}������k$�Q�A������ܩ�$n<|���
l���3�R�K�.�@:a���%�F����n�9��75YZZJ/u�J6�,�PTS3�ō�����L���з�ii�l_*���Ƭy&��h�d���I����<�נ�jwo�[H�D8�;�~��K&JD�Ν;R���j�F.���x��F��s�>�N3+)*�j~o��x=L�Կ$�C�\]�殜\�m�������z�I�y���!�֗�0�س��^��@��F����
����]�2���܃��r=>Rq����̡�������C�=9�g���<h0,��j6�_���ryZh�T����l��H���jzw3)m0���cR�^�
�#�x���?(��c0^(9#�V�����P�&�������9����.�^|#dvk�G;|�����?,��r��K���$�X��͸��ı�i�~I�7n�3:3�]��~��[�áQ\�u�p�}O�|�ΝW�!qk3]a~�?~�<���#q��$�.<�D0�����T�繞�FK�*� +�|�J"��o�(�H=1DLIE�~�1��:�P�l��+�[��8p��T���h����G�W�3^4�#x��YS�Ы�����[k�%t��Al��iOVbi孟>�G�;�Ȏ�z�C��2���͉�.pv�����vS��s�.���Zmsl�.�g@e~���oQ#y�B��4��C;��D*�(�E���!$d�E�?IgBogci�5�]��鵑�V#U!AS�#��J�#�����J�ZԐ$m4A-�@A�-�X�k/�ˉ��<v2�q��� y=M��c� wp������DUs�F�O���NLL�wgϣ�o`U-�/y��{s�qz�}�%.�_v
E�7h�&s�B��J~���A׸c'/Or�oދ�nmmͱ�SG��4�^4�@Q�}Q8�z.E9���ʥ�i��:u���ԵI�>ϓ^��!Q*Ϙ���{e[��$/�w@� G����F�����J�'���(/�6T�>��75� ��S���M�BР��@RY����U��{io�B�ܽ`v�'���k&
�.��q�&У�"�&'ZA���
::s)��=��/�#�(�c�C%[�kE�mW	�����˒�~�/Z�����Pq�g�u=�A�>�1ϘXr���9MD�:�(*C��`?��xQ"H��cAAAVOC6U=W
�*C==����?�ܵ�K�ҹ��М���쑯}s`�߿�r(��@AW7Fܗ�9@,�(�X��1=��0����sXSpQ��G~��zi���Ʉ]����T�E��'PY]�N��(ϵ�u��mU-�˪en���h�`N#�����������˗5S��||�7o���K�X��ӣ�$�@aqw�S7\D�f�>Jd.3/��j���2����hJr���J�N��k,�%T�)i�]��~v�-T�ɏ�'��[ ?H��g��o������:M@M�|�y=!�J��x��T��3�Q6��p�۵��&�k���&�N`!��]�b'`=��)�(+H����}�������Yp��A���|E��;'	��
߆7.�m*�X�{[��[/ʞ?ޔ�-����"Ք�y/D�<U^=�_���.2�N�5��W������EK�s&!!���ᷯ_߿{�f�hr���&%%ErmrJ���|��5�>%6����>�y�s�PO?m��P4��/h�f&�]�n�p.^!��� H綡`����ի9P8Ǒ�;���E�jv�{`�L�Z��K*��J
�����m��.�C��l���R2J��n��<<���2�zd���:�(�>��#H@�q�ę�B�EWxxV�	�-9*ji=�������fm߶�JX|�С��{��xn�.e=��.�	7�q�Մ��qbe�����䅯$�r�p���jߙ��f6���4@���}�N�,�����*�������ՓѪvЭ�� HH���L�3��\�|꧑��ngj��AK �Sm�TUNc�ɀ̭�8_i�C�$b�(9:�T��Vյ�HW���յ��9�/rX0 O�H���yii�ظ89�-���� ]*��S�
�Et��r��NNuuu�;V��Н��T��:`K�D7��'�N��_af�����������$���i`Ev��}O��J��U���M�z�8�|�R+������?�`�Tmb����y���O��y"�P@���=���q�^kW����ȭ����Z{3-�!`l�� 6��0
���ϾH���Ť%�r��EZ���L��I�SK�G�~Q��P~i+�jq��<F��m�Ӓ���.���n}�����:k�w��K��h���9A$XYYY�@�üt� �� �7u�-e�f�V�	f|uVRR:�sS��$瀼i���YT�ǎ#�s�i~�F�Wto�E8�/aw�*åKW�����s>�̱�A*��`H���M5��iE�vV�˟��U]N�x��Kn���W�ѣ�_�~9>4?7^IHL��311��Xn#���Ҋ�e�!ۑ>�ټ�|U�"zs����&G|E;�sD3F:ޚ��Z�\�㷎�N�
s[/�2��nٖ��q/	b�HLMM=�t�%N"�3�� 
��7��W'!�E4��\��:-%`�vM��ׯu55�G䍍��ы�nť�6L��W#YO�8p*!>ŵ��i)��a��J)ʐ�/}IO�_U2!"����q5+�f���n&�4�@�l�����fuBt�g�Xd*̢����W�����~x�(x'�_��)�le{#�W,a�e"��P1�>q�i�E�i����C�~�CCC�����T�~ǯ׈�\�rWRRRJRR�����ve��<�����H ���ji���*q�m;����X8��营!36�磣z�������s�����an�9�5K�����,R��|�ʞ��3ok�@Ґ�6��Ӽo�@l���].�d�V��1�'Ca}��gD�_�m=�]��-v�����}Sg�p�։'��䂫GZ`�@�Eh�,o �i�	2�a���/O�/�I���*8S�_.���b֚��J�s,q�����?9�=S3fm������40@?��	�e'|K�}�w� q���OM#KF�[k[�)9�S�QBw�W��3>}Dp�j����g�������Af��T��?PP�(�3-�dOav�Խ""�����-�H�����6��������I����h@}+_D�1<5/����e����Z]N!�.�/0i�N��u��I��L��!|vQ�}o%��3��_�E	�I&`���=0�hɒ��"�"���M'={�ғw�~[	YPdd:�B�x�DC��F�ְ��Iroޓ��8�� /��
�
N��0�)@.��^	@����Ȕg:�:PW�z��>od�k't�i\G��:P⢤���N�"�֡�k7����Ғ���ƻ�#8�9װ��)r"��	��<��Q���y�J:�c6X�%�E&��t���+���,f�ܷ�܀^�W�h~�׊vMd�O�Ҧ�=�L�dg��r��TI\��^�����\�^HKރ#���k�#�5n�/��J2��[��K�(ݒ""��y�&�a�I�}{LG����ߚ����;��:ۓ-SK�z�h��)�w���t�Q�)��"{��\�rC��M��`��ЕJ����,���l칡|Mv��6��������߿����ݻ�����%�_YE>)<i�hru��@C���9���W�˗/�,,m*:O+_\>1F�)~��J�h��� z�1�����������R�r�zp�t��DS�Lmc]]+����f�'��H�YBJ6�JGA��W#k��gG6�	m�B��<;Ƽ~����w{}�[d�LG�C��\�]�������"�E��A��G��_?Uu��^�	���D�u���0�V��eJ(�� !�:[����0�G��o��QIЌ{h��vGǐ!L�D��m2����!�~,����R���[(?Em�t�ҍ[����a�::��g���YT�����'�?}�B��O�r���8{H��K{�:�ŋb [�ȶ�v�- p�����7Z	����ʆ�����;z�;e� ��"��{r�Y�j=-���rZ�w��	II)`���h����%'WY��u$ܣ���7�J�T�J9!�g�9Xb#[es�t���d����A�<��FO��U Q{�4�_��^�[}��}7aL�c*O�\��w�w����8IFV��W�жA��m=�˔�o^=��G�>;,��6�wJ���FC��c�@�6קyRY|�!:�
��/�{���X��l>���Gx��X"E������Q�+.6r(q~�L�Yf���55����s�l
Kz�-�W����E�Cq0���$b`�P�=���!ܚ�<��1C��g���8p�Z� ���@�[��2�o߽k+vZ�����߰
�fҖ(���=61�"�%�Z�Ձ���qE,h�Zj�$jz��(�t��n���lR\�"�'�����klT���-X&�I�����77gg�OAye5�<����t��%�kW����͏អ���T�~�V�|�x��a� �Z?G�|mH-��&)P�~E�vvs�J`�U��>����!��"ӡ�g���B�C�]]������R��/����vR-�v�y�,��7ڀɰY��G�5q�='%-̓�\�!� "l��SV��9JL�@Y���C8����?gx�>x�P?~<Sz7J�=���LD�1F�>�R���2h�|"u����,��2�A�SϷ�aB�����������CY3/���6��`�@FG������'���9�C������XQII_j t%�GI;~a �rJ��d033K�N�a3�mld�����IMe}O+�=�;�p	�- ��7ys/1"�6f�E�g?���׺T&��\qo�P5�K�~LK�� $��en%Lj��d�qQ����hT�jd4|�,ʟ����5j�����	�o�,מk���Mf0����K\�2�8�%��Y�AvO@H�`du<uU���Tp%�k �"�~�]&@��z`+���x�J<�L�(��Bq!O���Wh�`v��@F6� ��P��v ����㜖^��e[�.��xz"8s��OU����s��
�~R��:�ߜdL�̞���삁U�ˀ�09�y��x�kp���e�Iz6�Ǐ�0
�A��^)0��ǎ}-$c�QN��x����#���� ����HA��=�B@x�_ݴ �J98D�f��p�L�Y�'>q�m��HTw��Nh+��ŋ2����������ڧ��!��X1��lmk�5i��'D�yd~�,X?����
��zv���&[��h�z��Qqy`~�+��5d=�Y�$Y�ǟ�Y(�Yt�? ��V~��O��g�ނ������s�v��H��)�9y��я����V�d;ʻ�A`�FO�x_���P�7w���7����I��
�������dK��������>�w2꫷!��3C�!�{��&׳y��;t��a#gh���d��� �T�
T�Ϋ���Vd���U�v�`��M���8�Oc�e�0���9F��H��~���p�|���_$ �cN\�t��u�MT��_,8\fa�"�h�3�M�)�= ��[��`RC�����,����FJ0�M���壶q����6�4�8:�[[[�c-t�e}��ҫ٪@sz��ؒ����k�«Sm�`�ύ����>�^f�u���{������J��q�0��������ߪ���I���f����G�y�=�iU V�uݰ�{phO��ޠn�P�;米�����ʨ����%U�+a��
jHk~:UI���P�I¦]��\���>H3�Q���-�G���k^��4�zpR�l���,��ϿM�C�j_˾G������1�e7�ͥ��^8yA�}w��2v���1��B�j�x��� �n�2W���`���	��w3���G�C@@r�h�l�2��<�_P�X��qo�#�5����-�b��	�Ǐ�-9Jמu+.��z��|Q�S���Dә�z�(��l:��e`8�H�_aJ��� �YX���͛dBBj���-J7�=�ՓR���G�gB3VZ$���7^��F�"Ga�O�ѥ���l?|��q����	>�=6:��14����g����X�Jݰ���Fý��oN&��eT���"���<����T��^������P�% <�o}}�2u+�!g�%X��L�Q˭
OR��%L��D���/ᖡ� ���Ǿ!A�!��]��.&����8C��"h� 4��K5ݛ����oy�ud�"L��&��b<XZ�I�(�3n���L��)z~ j��4�$�c0 53��M3���P���������P�:uJ��E���ϟ᳌S	w٠8`�g�Duc�jZD�����̱)@݅�޲��N'ğ!�.qFҜճ1C���B�
E��`���7翼��\��_���~y�?c���[��#G�(����$�RS3mI���@7�`^ �������t)��̯�g��_�-pJ�����b%�~�C�A;H�v�1��<<ɾ�t*��0c�],Im�v�c�Ev�C���rssMMM�oȿ��B�p�g��F�����N��� ;²� ��o�+\��w�_�4���?���3���}���w��%v������ٷ8��t,W��4-������ū������L}��(L�}�w�O�kega/�����Yq��DD�8�IFY$=(-*�HB�+ڡtH��.wP����hjbR73=-���A���I�%%EPQE�� "��Okjɱ�S�u���G�����P��mY�y���R��'�S�ґÇ+���>EGG���8AGC3k]��}N����}0�(�;̍Am\E�Ӏχ�?{�'��Wr����2]jz����Bv\a�V����df.ܶ��v���������>n�ޅѫ�e`�61_3}���ZhP�X+:�U����{��x��4�9,S�i��%�}�E��?�:9���#{w��m���w�h]b$~/�1hdmaP%2�cG͹�]�����W���K���FQǔ�[��ڴ�;��t��0n�^���q��X������?�����ѝ���F�o U�\��@#�L�.��M2��ȼ��sn�z���+ܱI]}�o8�Ӕ��P_��n�0����qs�%;��c~מ�[y��c��d�i��\�Jܾ�s��uw�}}l_H�\�d�t�Ѓ�'��W9C;��f����3���le��L2�,� ��;���ԧ�D�C�Â��2�x���w;2��d�[{��,F�����;���ܼ�yw�nTέ4�,`5!�^��Spp������)�� �B�t�@14�Mӡ�!H������-$s;D���b��ݷ:`�������,�F��m����{��X�^���� v�Xv���w�ky�穋�R))*��,��� ?J�4p7_ad���3�U���o�B���M��Oה�� ۽o�+��V�(vٷ��-A��_##e��^�Tժ� (����>IKN�R���������!Ӡ1�_���ST�c-���?΃�c�*Y����\Ft���c�o�!F�*�#.]�G:	�тদ��. ����6��(���n��1����wo��n�����%&%������z�U����ӮÔ�� l�
����A�cA�����stt���Y7g����b��cs���Q���֡��w��W8j�޲�.x�2�l��ژx��eMII��ty�+)��<������� ����uzxj�ӥJ�(�.�W�������v{�7���F�a�E&�"B���,%�_�~}"���/��8�mf�u�{:�ï���/��d�)����)����/�����w����Ą\�5��Էo��A\tq,X�4�39����������J��X<�V�Б�=W���PX�Aו��n�τ��Lw���ef�
��ʆ�Ye�T�-//��φzROqqz���!l���P�7�ͱ\���<�~���|��MZ���Z�I��U�ߙMK� ��7�tf9�D�PQQ��F�y5���5p�7�e	L���VŬ;s�F҆�1���D�6����J}@�%�(?2^΋�vjXpрN&�f��݁?6���3G;��j����
ZA	f�:1f]�������o5:v�����Ԕ��5;�����Ҡ����o��ٜB��+W�|�$�u���/e�U�%z��������uy�  @V�C��C�!�:���"���>���-JM5���LS�P��\����olYZ�j|<���%:�VH)���~ѿq�m���U%�>��4��9�W9
�۳�Y=g�y�>q9�4^_�FD����\�͛ϴ��.����P���r_c%'	Z�CסTY="/))9�4R}�p��>@�h�+c?)������q0����4���5ݻ�����*b�v�,��٪�ie.�B��+�3�vA�.�9.�S,c����z�������傘�1�߼ys�R�����������8w���K@k��>��������*[�0�)z�t�Dlssen(S�[�f(��q���L�H�'�jZ�Ipo?!��"�Uo��E.JĤ//:������z��T���#͑.��~wC��S�+KY]]=!..nm��|WN.g޵�P�\��E��r	�ݭ7Ër`��f���j4��[]̸͓�`Q����(�/p钞��٬p({J��٤�/h�me�Q�q1/u�`Ӌ��r��Z�jkkѱ� v-t��K!����&ehR\���
t�g]φ?�)S~�b�4��rɰ�9���փ��s
�Ωc�q����/����S*���u�ʕ׏q�bK�l֚>��7M�y&(ݕ�D�3C����	���6������;3t���pD�=�,D�:SH��������ѣG���v�<NL�
ڋ�Uh�,���KIY9��iWz 5�t�#�-;�|Ok��?��>��(�r/>op\B��?{�<��{��0�в������}%-��]�v3o��_, v�l�	���p������|y��]Ni9�z�??�hҕ��I�j�N@pp��놯��>7�(ZU���L?�G�#��m�f��A-]����N�`Q�3H�=�:��;�4��>8f����99��^���,���� ߃a�P�N@(j6\��8IC�V�t������e�6�fZd�	P0x��$o��'mT`����\���GF!캅2ڔ�;D,aV�cll����ԗ��E$3�E�G�^����D���TR0?+3�>[����[��פ�0[�͘yO�����'իX'��חB�ļl�^!�2/���]��O��δɉ�am�Z/U͕��
�X蟮�t�����S�/����3����qp�FP�����z�c]``^~ND���@~IIA�[^��P���� Ad��5�k<]����,��)@}��z��	����10e�9Œ���� &���/ {ĝ��X&'�� ڍrv�DO����nՔ�t�����;��� ����g��l�p��ú��j�.@���DS���0�I/ "�����1����ƺ(ZI���mc8~h7���A���!�"��r�����&�����y��H��b��V���L�^��5���.1�l*^�E�7��NC��z{����������uttD�ʲ�3������+;<w�f޿�@���
�d:�!8���F:��'z�������瑂(���@�S%���*زO�C/ȫ�u�����7���-x�;(�⪙!��|O+b0?�@�߾{'S+u�^>�7W6F|g@ yX��e�y*���g�(~����U�VR�0�ֶ�DS�\��r���k�dŭ ���J����3���JBCϤ��%��tN�%ɕ���P�WVW��{@��-|�E�KA�6Ʌo���a�C�Б���� W�����y��}YY(>�B������ֶ��ly{��-�1%����e��EkP�鎔`<�tI*�/�t�WfTc��e!n�@Nf�n.G�wөFB�pD9O��Z���Y�n����1��=I�v洶xD�o���c�
-%� �v�����p$~�<ɕ�]. >n��@����$ڞQQS������-��M�ݓ�����G���G�/|~m�dY�Ul'�%m/�3��P����g�^����e��������A�p��Z���fҷ~K\�[��t)Qi����1Y�Jq�!\��jjЋ\��j=��R�ٹО���,����t�^��O��S�G��	7�=�e/ѝo�knk):� B���<��ě�������;ZZ�a(�mp��;;;���MZ	D"���Z�911Q�H��G�T�u�8����$kZ~;�%eR���C�<�w� ��U���C+��+�I��6����}��'%9�W������#�^�|�$	��r�'$T~�E�b�n���g9�B��1k�Κ��@gy�ؠ��"��������^��4l7��OL���W,"��J]7?�7����-�&|�q�nZq�;��CЙADD�	��ݻ?e��{�^�g{l:��M�v����/���SNU�z2X�4j��h�$~tt�uI
�>g0�Y�cR�Esy}� �gڟy���\%�C����;2�@ȱaBNY�ߏ�R֍,���ݻ�A���ж=�"��\`Ɣ���� �M������Q�m�/a�U!�6D
k<x� G�w��+p�o��뛛�U��:�,���ղ�&�);�D�7ߠ�8n���(�'G r�d�����u�2XpV���������f�^g�Z�=o
��g���(�	}D���*�9o��į��͑��]i�,<<�7wM��P.|B��0���Z�i�7�A��EcQ��z���z�/�"�TR�xAD��{���P�������޳�w�^�I�q7�	B3T�_9��W���#U���`��*�?[�Q�B��H�L�󭬷�g��6
ϋy�@���:+R�3�iݦ���d��;e�^�LCVMY��龿'!( p�s��Y
�"��^&�W05�Smǯ�������<�|{2\�0͞<�q�6(M�믗������m��GO2�z�k\�|���R�kJ���^4���L�6�_nm9�噅���nT��%R��m��_�_(^�t횲`��[翤��+��V[�v�?[gg��hN����*���� U�o޼�&� p����1g2���� ����j�C�+�����x�1��~��붒�����6_>�ݮ ���:V��M �,�	Y�NH^�o�9s��LЀڢ�R�uyy�G�>��� {�� 2�~�����B@/!��Ͳ}�N�����C:l����?e_T�f�}�őڂ�H� Бg��њ�Wmƥ���4Rv���Z�7{��sB�d��5�u����0����$QDz3�ٗ.^�T��:U�c�����f���|��[��?/Vc��;���*W��\�5hǫF��-�x9۰9hu�v.�������1�Yp�`f�S`�r�F�t�d�w����4������n��<F@eY���{�nD2���P=:66f�=wut|\DM]��y�Xr�����z�`º<�OS"r� ҳר�J�X�`�7�rVNS��v�����q���ύx��v}�^�ݺ��#�޾=��Y�����#st/�wƯ�"��� �EDD����㱟U埊���f�%pp���4
�6�U�ް��EF÷���,�_�d���T\\�{/��V������\�-�G�bB�%�I
a0KF,��=S��Yщ"���LvE������l�N��}�D���?�����ã#Z2�᫾�N�����)��20o?�e}^���T��mwj�_.��q���ꙓ^↑N�$���q�<<<9� ��EQ��sYiZE��@�M���L������LI��T������x��w�@�́�RC4�x5��-1d��c�pc?M��5���0Ғp!=��A!���|��OMc#��E�����nO��..//���5\R�h࿿��pm��z�p~#�e=:�ʽ%�H�(��������a����Eyyy�ʐr�ED��m����)���e����[�VUpr*H��6e����)�p�>G����G����0��>�]澟fڙZPg�%�u�����iPL;�:kR����X�Ms `a�ԽG���\Gs�dۚ&)�ݸFtE%U�ꖮ�n�=���lR�}O��H���#+���jٗ����� �����!���m,�l'�߲�kn�b:��	�1L4ci�1?��`��TH�Q�|��X�~pŰj�as������\����C���\n�7��~W�f2]��ZZN���C4ő��ݠ��!�]��\�LA��5�h���z� ��+ͱ��)	��_Y;L����8wL��[����VɫBb��0����2��v�WR��~�ldkn>/;wz��ԩS����:�_��E�q��U����r�M��az�Q����4��$+-%|h�����-�ZE�_�PPR�K���xٿk�י��K�^6�D� n�3���+��c&���� ����p�Ϋp�@�`hjH���ѻVVK[^�﫪v'�mg:�d��V�����b����L���WW�*K��;3�9�s$JJJ��ܦm�2�N��߃ۦ\�@0��R��7D#�>�X�#�O��c����ģ�>��8��w���E F ���)�O�5�@k_����{P�V�r-�//߂�)�Lc�� �x*��*S q�N-�D�ů_��2}�ԛ���}$b �Lll��YY���9�8�����0-II�����`T� |��?��F[$�)��;����8&"]����Ҧk���cG^x�:�'�R�h�"�xT���r����VVV������0���<DW��N_L���1N�H�Х&ɗ�"ă��ٕ�����PbP��q���������Jl����J���j����:�N����L[���{WJ����YiN��.�\a��,��`$����/00!B�sU��Ý;��^K���-s������%��&N\m#箛��=�mkJ7�]����`����}ѹ��w���;��[���$Q&,񀧦Z~Y���vg�.�����!�OȻ���U��-1�	Y٠��O�l�/�LDL���z%-��aK��!*���.���G�9W+�a�y��^��j���
ڧҸ�~���ى2Kw�]4�5%$_��+�IT�?N��a��Ĳ���-Cv>�7 x�ȿ#��(�e�r�k���0�.HӺ�Q�G�L���ₕ�^���6�'i�$^��~2 ��%4�ŜK�յ8ܮS￥������i���96?X�^1\�fN��u|��bt��J��N��k_�.Yh����dN+��I���k3��X�?��)ם�j���xA.r����0�j��:���#������t�Y<�>�I�:9x���fQ���ߏ1~:C8��E��~/��f�-��6�ϸC$/A�'�X���020��=��`n���W���$؂���珐�[�9�������M�/�
=B��ڂ$&���S0ؔ���$h?������y��m.?44����8�(-��\n�w0��rj^� {����ز����b�r4<��L`��":_�hܣ�K#�^�N�0o�:D����h�̻���	��vqw����Z�R���1|�h�&��#F�k �nV��k7'8�g� -)�
D����[?���j���?�|��\N[7ɰ}�S"2�Oc�FX�@f
ػ�g��w�Ɇ�V�?~�02����{V�=_�����H�l��O�_\� \-�Z~MB'ԍ�e�sY&3{)v��R�:�\A)�j>��3��1��<�`t�;BW
5�MNT���5�C@R��O�r��2��� ~����P���8B�^�GM{��7��b�uMMA�(��?�h6<��\�v&K�ٹ�U5���s�MNO�U��0Ud@��)*Q8�+��������8�n����]�
ۍv������Y�ٹ�>�]3�ʊ���N+��wM}�zۼk�U������U�nN|B9��˛e��\�&�>:1Q�o5B�q�|��߿�ҫ���Spgels"*x�Wt �� �yy|�F?�w���67�Y�Z�1�`�����ҿ|aR��7���§�6�r�[?��<+E1Q͔����ׯ���}1(v���s+l��&��7Bb/Y���8G:���$H��*�QA �6�:h�Q���Z��DG��@�<��&l0��Nˣ��f_!_�M4E�`	u>���Z��,���v��I��N�XC��j&^���������c�s�#U��:�	�ppX��r>󰯓�`����Zp��dt�v�.---��׀���+8�G�}E��f��mms��gҲ��.���]E�h8�ϯ�W�vS�����>�n�f�II�Ů���"��[vW�Ο�)X�Ce�A�ߪ�ؐ&Z�$��q��k���	>EI�A����cQ8X.���d���k�7v7
�<�A����:r�Z��Rm�TUݍB�[?��i�r�����n�΄l�DBii���p�?�P��0g
$�k��v`��4�ƌ~TW�3%Y�yrpэ�]Y�s��)bI�`Mq�To��k�����≍��,��-9���S��ILJ���D�Cy���w*�Nw�_��蒑���n�[�#����K�m�m_%o)���Cf�s����g��={{{���l9�kkj~6q>�_���m�!�� #�đ9�r)�qwj1G�h�țVPY����^���k�9eTsR��^�咯���,�4	jL
���g+E�ϋ��'�i|�ar��
J```�k��{:O����;šJ��HH���H=y�䎸xUA/����J���АE=R����g�YV#�sX%Z>So�,��`B���U`�r۷DP�@)����b ea'�	͞�g/����ROSY�?FS~�<�j�ǋ��`��(�h`X�YYg-4�4�Յzٞ�]��u?�������Z������ 6Ts�#~BҎ^��k��`)
�d���-��S������w �܊ �D0�cxћ����~�«�;�F
����ͅ���#�frg��`�.��h����	�W�)�8kr�����Y�"��S�tŴ�e}}}���F�h����l�{��(�U%k�,鐫w�(�u����ga������@2u�%
���9#'g�|��G�5��>�H5���s��z��-����}�F(���K<�@3���V,��廇�|)����Eq��!�c3�^�	F+J�"h3҆�&,W���%_PPp�E��d���eIu�Ѓ	@R쁼|L�W���Uq�e}U����l�������O���Eh�"<�V✋--����� ,���#�'�:'��-�zyz[#4F��7��jj�3!k��q�w��t��ud�Q�%�Σ����,��mfh�ze���L�bL�u�H�x�`޽{�&{��H�o�iF��|�d��t��b�F�0�����7��կ��\i&?��ٴϟ����y��64�ǉC�ހن��u��r�\?� ���sk�j��|��*���U�鉋�F0�?��hn��|ę��-z���(W��������8���ۨ��
�xD�k��r�5��bI���p�VD��t��>�7��لp6u�󔭶���g���  ,?g(��5��k�9W��t���5 ��.�����h\��D]v�YIɕ�s#�x�Yo��۲z����㓓���"� ��?"�eO�Y}�t]��խ��[�P�n�C/S����ٰ���?ޜ�0��5��_l}w<�o�����Rf
ɦ����2����ݱGˈ�dš���ǱJȖ������s�_������s��u}���~_�W�C��T�����r����w@]]���jǫ��'�P�^�zU��RSmՈ`�����]5���bb����?:�{���:Q)�]x�ߤ`ύ'�ѷ��E����{���MQ��-3��R�˅h����ʚ�S�#��E{�|o##����*��	�j{LL�����/��8z��lYf�i�ؗ�LĖۉl&zzCu�����9�k��PE�3�ˏ�ě�����1�7�J�D�'���P1���Zr���q3K�_�l3{#ZL��5�#�U�7����p�I��P��s1��n�����r4&�`QҞ����}���J5�!�-:�2�8N���;Q������ډ���iz�@��;b�ѷ��ĵ�p �;�bK�VrV,s��RZ��\�2�&I���=�t3�R}�yu81�P�U��1a7���=KbA�����q�d"����!�Oğ'�Q����N�M)^�ǹ�����\�ݺ	~��l���2M������`�5���ϯ8==}�̙���0������,�R��8��ɑR��E�i����ɶq�퟇PU!�t�`0<\%|��f��뭷��/����Rn7PM}�L��$y4��~��8?�����)��Ӄ�QW	�<��~�q���F�Ѭ�Q��h�0?�1��G�;���������e�v6ܷ?9W���
�<M��D�x|\�[7
g�E9�'8e�AѻTg3��΋+�s]Wq-�s���_|̷�'5�o���4.�@�%܅�oWёE ��o��y��ُq�BS��zz187� .� �xt�fg��ɱy��n].K�ZU�3�0h�l�܂����{!��۶@�����v/~B�G$|��莓Ԓ�,O]��T��'�� UUU5	�(�Ք�ɿi�[USs�����~a4�ald��Y&mk����H�A�D/��� ΀�{�w���FG�#��j#�C{��]EE=��t�9�S|�?�T�`�d$%��\c��/�%K���g����jH�s���T��ʿ<�c
��o��<	J��#g�'1L���Ǘ@R<�+��ۣ�:�vR�.���9;0��Q�dPL�@������'CCOݹ݊���,7E�̓ 
�	�t�/��';���U�
�\+m����1��� 0�[I�^Vf�mtB��Q���fI���x\fp^�hҕ-�-�̣q��a��}	����ܾ$$�gt��B�+���}�~��&IjK��O���]DV��e+���T����|����R��V��dh����
@���̢�TU��Y�N�?��M�"v����.7�1�;ުNX��	�z�u���vh��MKX��zb��T�ѻyꝧܴ���0@�Im��������@s;O�@Yw˅	8�B��5-#H>�N���(=~�d��x�
7Z��Rq���W��ޓ�d��I�
�L�����6�ZZ��J����ж�i(�Ҳ�޸*׼�����`ͷ���3�Zl/��sa0}��':�����|�����<T'����Ƅ�H�fg�M�U��/�s�u�v�\��/%a2�h�wo!,U���K�����N�����d6^��Y����="�hQ�81))�u����Z�J+F�e��D��R��z[5C�b�q�	�ޔ�y�1P���4���V�<����j�gPFg�)�C��~12���w���g��`�ǡ@�-^�o<�Q���`��-Ӟ*�ڳ3:;{��߼���y%%��Ô�#��������y`)�9989�6��Ov��><<<�������6������7��&�ѣY�h9�յ3���-O�4CZS35l�9�~Ag{Z����ל/�t�*0�nDfA�Ɇ�\�k(Z(��D���%���
`��:@of�m��iiw��
�y�@���A�h��|J��(C /������.ްis��)��6��j�`���l�2 ��>��S��Y��	�O���Op�3%_����3ȃ6x��Š4Ի6ic����)��0cׂ"��H���|��H��6�ѕ��vsZ.o~��O�J�,&U̐��$76>��쥤 ��.0p�ΏB��9Z�,��
s,�_J^>h�nk��X�R�>J��v5kml�����"�Z�Kx�����V���{���U/x(�Z(H)�L���/g�)�V�9����}0rc5 �V����+�qÇ���vӕ��u�$KܸQ�զ�bI��W|:~�<��b���L��!��
��kK1��w�^4���e���2 F�[|�ٱ'�F�"�+f���8d)J�궑�Af��u��d(p2O���{�r,X��Ҍ+�,D�r������gYXn���?S��s�q%5���)A��4Mb.A�'~���l�aܬ���c�8"Q�G))��P�x�n����?����<~��h�͵(-������a'^���.RAW� ��0|�/o<���$��e��1Y�0YM��v�4��t �������j��G���X111�n7�����bH�%���m�`a��b��Z-��ZZZV��#' N4@i��s�$_���w/�Z:zv�R�<��;)����h����;m�in~�[>X���)�"Opz:ߦ���T��0�')""B1���o�+��@��,,,�q=�==���UQ9/�!��tt����䦿�f�l�%�P?F����`h8���μ���!tFP݆�����ÊI$��~�B��ь_�E�FW�.�����ՕcƐ��R�*O~���W����� �,>��Bk���	YX̬w�P>5����
D���Zե&af��GV���!5+kN)���`^�6�B����lkd�AL� �X"�4��3��6`T0��S
�Z��"�j�����>��ǈ'�k����̪�����]]eS2�̬����=Ӷ�;��m~��'�O�а{zzn���<zt����������k�U�vN.���b�����?~��=�V�����:cRvvK�4�g�+�B� T���%oc}e�����-{�"x2��Pc�3�\�鑥�6�������8�[�4dQ��y}P������y NG�xzy�|�rÙ�-��n��M#X�:�a�&I7�-"��)>�i{m�
��Ž�s��v�X���G{t���cbc��_2F�F,2����$����:��hY/��ˬ��{�yfb���kc�EY��z!|]q��6�Ho:��=RP��|�NLf�]��yj���_Y���T�dF��G�"�&\j�ꊮb� ~�b��d\aDK��8ղ�d��z.UA���=�A?�^��!�_&�Ro���UCc����w�2op���W���6���`��ƌ���hP�_2	��N����-[�+�ٽ1�G{!����B2��~H�܁6פ��}����F��F���� }Y��k���������I2�_՚��Ϡs�EǄfC�H�.]ZS �L5��i����N��΃y~�Լ^ohd�(�μ��8Z`��q��hk{�oS���蛗.^T'�k�t���ǃ�_B	 7@��XH�b3����
wq�!|
��w�]tl�zʆʓ\Qjʪ��ム��s�0�����-�6.OT�'�F�<Zܺ���FRe���t�ƫD�6��Q8�]�s���`O�7G.�D�����**(����Ԡ��h?�]+~XB|��W�+@>�^�zE�>�������ղ�hj���6jsԔԙT��+!��`��Zk),�斖J9A�9�	�!�g<ԁ/���j_�ٳh~PޓZNN�roSU�n�	8`��}sN�u�$���9/ ����a����S�~����e~��'O�@1}
\E��:��u�0�xv�ӧO?�\�<�q
�S36NЋHL�e! ����O�"1P���5x���l��a���C�
�.�%�h�ϛ�ƻy�ƈ]t�iOAa���	^,�#�����Pd9�F��d�sƸ	jpMs�VJY�w���w\&�D����܊C�Cf����i8��	1W=������J��2!*(ǩS�6���Ѯta[&��{�<z!�p}$�f�2�u2	���]-�d�Q�BM��ty���ƞ�d�Q�IG�tSm��/�uh����{���B�F�Rd;�D��g4��Cq����ۯ�~�زH=1]��܁̣���W*�d*��6�@�2��B��W?�ĔE**��Kwf���{JJF�� ����S�T�lޤ�H���a����2�3�ˌi�̯`�M.^�T���a�	�8R܋F���T~��ſ|�Eq�`gI��ϯ��w屩WlTV��SO�B�
�Ɔ�y	���۷����Q�`�\��(c�:>t� 3G2����nNt{���g�p>���ie��R��ٔ�����C�~hKRV[U\��W�w����ԲM~ʧ�����;p��)Q��+!6�>|K-��$�4���p�C��{E�����ԧ�+����A��3:��������	[)��@��q���C`!��JH�2���J��ϫ嘶��xC��o*(F@Wt
5ut�!�eJ@\8�
�I�Mic�#d|�e��
������1���jNj9�AW0"jo�B'~�o ��ε �+)+/���1�����JC�W�յ���ڡ�[��A sM��94Y��BT���{��;�'z
�@klN&�NCE3�S�����[R�- VjG�	<%�e*�4x0�s|�?��5Y�f� �&(%��[���mX_TŤ>���E;��~�����(B{����;R�rccc���+��s�q��\��˲ 6o3���h::��8���������F ]\y~��M��:;��]��~����a�f�	4��@t��<��]i���fV�ښ�U_��8�7�%�$ ����ٕ+�SC��M�6��~�C�
Z+o�5_:aK�@d�5���(n���J�; &��(D{fMgn��'??�	@Hoz�M�ҳ��Pu�`/�K����A�Z�,� ���V�K��ŉ��^߷W�?~� �Ҿw�t���y���1_�Hc+�4S84�w�<iApr�S|�-��Hi9�78�b�A�)��2(lh����S��П�U�?;;��}+t<�"���
6��&����znn�;⛑��՜�"��3��b\�ZڴOR�w�����94b�%2�O��T1��H�yR�����P{�;���Tm6;0��ou{� 8��B���ء����ϟ��\z���72ϓ"���e+�E����/z�E�S��Dݼ��X���K+游D��-��B���@{�{w�"ǹ��6fm�[�ܡ	imD�x	��\�$d;/�[�7o��̇^t�`��X}�b�W:T���&#�D5677���\Ϋ�����lӰ�ɡ��Na����ϋo,����w"�b0L7�/�6\�l��|F�;Ӫm�F�^P�~d4��<�t^�/��.�����y�;����� ��?���dd�t��z�8��/��"eL�vv�G�M����a.4���8��K�:{��h�2�E��a�y�8�OE`�d�C:�rP_ܠS��i�p���x�����t��DD˼N�0�v����`�����@\J������Kˣ�8�ص�y�	���Jw$������Q`��L@;�YT�Q�nV�S<���\BZ�A�5�����	Hױ}��J�.�v9Z��h�؝���eq$�"�M�4Z���H�C
����`��$1}e��YYYfO��Y��d����[�~"����70)�K��-��N9�-ii�X���[��V��*FR־3�P���c��8�0�8hҤa
2� ��vW�0it�Z�����b�P������l�����ݝI�����Fe�v��|4�{+�0�c�^���C�^���̌�`>!������b�!���=���eB��ݻ�#���M:��}i�<C����f����+��P3s�����)�oK��\���_�/.&�¿�OP��o�<y���8S���N��zS]���j}���ҹG[��MC$)�?�.Zm�-�5�~c�W��-��U6��ɓ���7���b��P�Z����;���F*廎��O:3Go@Ē��[m�W,E��:k�|��1b�W���B�E�f��^Nw�p^��]gA���4�oA�������Jܒ�?A�0?�e�&�������������n���̌��늁�h���˨����������� �9
�@ȼG!�$$�mR�G�~����H+ �<����+j�U�,��
�A*���׃y#��:S���M	$�[rr-�5( �6��8��HMʾ�x���`?�AG�43��l����T����[�0K��Uү}�wsske��er�!��n�zT~�����&MB�p����}	�Y�.��`٤e������TyII��4�|���gɇ��dx�L�?�����e�I_u�P���3O�>ʭqi�|�s��'�~�Z�2���z'�,C5ndfV�;2���ۛrs�N�enػZ� �1��tim]��j��E���o$�$˴�[���Q�^=d_a�c��Z� �	�VEi�bKP������S�F�F�eځ������ƚUTTcs���.7`��u�v������'(((.���۾��d�_�w���$5�b>�}��gGr��F{���(2�0�ٛ�@[��_�^:\&�0��P�g>���iI��f���]	�ޠ)�jttt��t*�m0M�͙�S����F�mi�U*�4:Yr�hdb�(t.`!�&? $�<:���^f��___d��Y��t� ��;q����M�L 4��'۪���I@��b�f���60��X?����Dl8�$��L�&��uP.���@o�<x�Gl����l[���(������<w|fzz�7d.�ilh����už��R��Y���u�������ŗ�#��[���G�"����۠�X�(c�Ƃ���r�?���I�D��(���h �������������P�V�I0�SjS��jhf�r�/|QPP<�?C��f$� �D���0�*&���>))��H�ڝnۋk*�ќD7�s��K�M �j��N��$m͝�X �eo�t����R��d]������ǿ~�3��nf����{��h�9�4��.�ۤ�S��w%�/�����M���MB�[���u��񺴭����pA�� Gh3Cggg�
ZW|᷂.z���!��?EBJ�X�i�J���˄3�ݤ����m��-.���S�,"b_�;u��,,�
�/�����Q�X�"�W��qe�
���l�8�u0̑#[s�\ڷ˒::�k�M=
	ğt����r�.]��HGhYs>p5&��� <~�y��^�2fN����mi����3�k-X���������hi^P��(���Ԑ���M	A� ����n��ډZ�@*Z����#�`�WK�^0��̸��63r�s�6��kK3;!��Eu0������9d�x��T��l��û���C����hi�@l�ˈ4��L7���&$o����ɟ�����4 z��� yk���8������Q�D��
�j�����r�ᇯ��Ê��4��@�N��J�|����F�prr� �iYYY��]WN4���R���ԏ
R�b�f�?C�>"kd�r�O��Bz5R��A�*S�5�CrK��/mi����W��:��x	�'��ހ@�}`���#�����ؾ'h�Κ)��i߄Oni��;ԩ��r�t��3t�n�J��h^[&��T�y:��d�ӧO�'��d��b5�Q�~����yJc��o���إ̬,�dbC T�M�Ep��5Y��%��UT�a��?A��vnm�C>T��ߊe�ֆ�ñ��I�$Xmmn��(���J������J���Zi��~d��W�@��JB��޳s=��5<��N����� �S�Vd(����}��ɜ)��[`�K�4��b���ğ�3�Tf�d\G�<�� Q*�m�N��[�nQ��%������==�*`��h�BMM-<P�ܳvR�d�P�FƁ�7]�""X���KX��r��֖��v�����C=H��$���r>q�p~�,�J�?Ґ�V���.jho{��_he�y�ٴl|�|x<#Ҧ�5d2ϊ_L�@�;ƾ���"ߚ!�h��3���u��߂$"��tV�����@�a(Hϐ�_r�j*��
���Cp��V����ȳ�0p�9��q==��p�1�{_]�X�Ǜ�2�_n����+���l{��9�m�	�P:�oE����YɃ�_U |`�:L�̪֘7�����c$r>}�-���up��k�r ���c]5�D�>> QQQe���摏�w/nv&d��:#�a��;F@��O�^N,�]YZ���e�z��$y����ܱ}N_����M1d���[��A}��Y��@���V0K��H/7�d11�����������C�,�������̐u��$�eR����ʲ������4��m���ў���m�I@�:���:�@
2�P�LKK�Y�T�4I�Ίz�f����W�[O[08:\�5�'[����B�Н'�I0��v%�e�+�:��Ob�322��_�!t}����u��FU�ƻ�A���l0���/�I�^j��{ޡX��¨��.��b��֬_���Ɖ�S=�`�x�:���\w�����Z�+V�&~�b(�C�<E�U*�+�~��>"q�=;�gW��P�l���.<�/���If��ϐ�D�;e����ͷ�f�D��߹�F1��ˋ�=��G��1yl7�`i�Y�w׷������Α�?��~jBF�m���qc4�^��O�y.T�>�SW����h������F�o��Ta�P����oo�}%�~>&��z�7e&d2X+oYZZ��E�zF&l~f?c/F���_=��6���S�<�G��
bBCC3�p+�]C�r���=����@��7$G/��`�8*)�k��ڶu�d�\�!;D�% ,8���g�*� �g:g�'a�NhY�X�l\S���)�,=�P�[G�P�6�PSq��F�����"�QJt>�|�ZLO�A�}�p<`Okl��Μ1ϖo^�N��y6�S��ꭷ{R ��k��S��k��g��kE�M����s�Dmu������Qki�K���N��3nڏj*;S�	��q��ʺ�&O�e�}FhI��5�:�)vSY>Ǻ6=:�}c"-,�Y;(c��gi_H#�qP�[�/���J|4Wx�%��F����NQ�-9�L��-gާ���^ յ2�@iU��}%��M�;��8������;�P��D���D��V��o�JT�o�F>��?���^m�p��G<O��Hm	]�!�\Scۑ���|u��<k":�c�i�+�i�PI䃵����ᬂ�釟[w6�>s8��x3R���D�0Y��m�꧘X�OY�*Fe��D�A�0�dU��ɗ]�:$4�b��h��f![�����=�M;��=����/��Թ�˹|xy��Y=L�����$�[���^c!�<�$F~?kn�z���~s!�e>�q�����:s��p�y��'s㩛qSLS{��Rm�p7t��y�߿�9p/�&S�l͜�Tz��<e�>��09u�+K��_����~������T7m���h��-t(SW���}�:/�!�$���i���B�Ģ6s!Z��-�8��˗���9�n!D{�I��-��mڲ���;&��6ފL/''G\��ئ�x��������!��CPe��
�nd�e�����?z#HC�[񳻻&���-4"BS�:������b��2P��mc֚�Q�����(B$�>n�+}}�̣=oK���������k�"e�0��k��?g���$ւ�D�|rK5y4W{��_%�,�������3_B��8����@��@N��SF������Ҿϭ�!oZl�S�J��n�
f����A[@���6�.��\��g�����^z���o�E֧��#޿�C3�-��W�q43�.۶y+�p���{��#|�m��yA��������83C���{�i�5T�����䝣;g�n[��؀c�B��3�1��-�\�T@h����4�Uj�"O=��>�#�T�r�p��M���sn*�eJ���Ȃ@�BZI\>nf�f����4)6..먾�ܳ�q(�v�2Ҧ?v�T�w����}KT�
������n2�mn~�?���lz=��mEEŒ��,�>��p<�������!�	'�L�Yo0*yINV��64x.�G�f���X�+d7f)u}j7\��\Ӵ u��g�]*N��8�1z�o�k3R
�%����4�=��_��j��<�����yV�����~�[3�ڂBQ�}X�G��	:��fQ�Cb�Hn�C��P��UO��WQ�m:`�4Y���G�.Mr��������Q��O	�V�����e�㮵�*�V��@�F�)�0��縩��A?����Yn�)!�l`���/��c���buԡŵ����_�GƦ����օ6��n&�9���\58��w��Yo��&b`+���������4	Z6Z�����+���� �w(���Wj��\�u��N�������C����{������sԹj/[��:��@��C��t��#��*���pm��1�-�C\��0���쑉�?KF�L4Q�0����>�������4% "re"���d�?����MC�D�A���H�v�#?߃&��{��o;���)�?�fq/���>{���)?a�P�*����Ä13T�^q5@�Og���H1 �zt
���9��MD�A�'C�x�%�mҺ1��ϟ?@��1%�h]�zUbO��g] �A۽"	<{eL�Fs0;������AA>�O@��652�W =�����ɐ�6�o�E8Q����!�mlj�;v�D��M����=��h�<�s7|���͔�����J��=Z�nV��/�h���AO�fgէ���=�����_|��8*���v�xf��`[J�3J��������������������Q)mo�n2$y����qS^%}���@�_[uX�'^>#�j׶]XGٛZy�t�VbkW�]�;EC�Tr��ٹ�� ��P�&��d@;y�OG��f�	����bZ�.	
:�&~lSS~QN�Hek�t����^�
�DV˄� wo�����N���xy�l�lFU}�!t��Yq		���:�,��7 Q�u[�Zr����{����Wr��@vO�m�NF�g�2�5�<� �74��s;w<�@�gn��݃):�GRB���P�9�4��$ pݪ�Ot���M�Q�����Dw���x�K*[�K�O@��S���HG{�m!�K��Ši�?e�xP;O��O�\\��z^�(:L:3ohkk+t�p�b�1,4��Kνw��3������'�?{FFz�����3*�ުyDS{{{��q�<�H~Jc�W���wYXY�/��Q�0�1�z��
fڃ�qD����+����u�*|�jب)MQx�?΂�X���o~$��C�}ra�"Y�it��ׇIDޓ��ah̏�~��ݻ���Û�)L�,��Ϧ�{�l���'x� Y��G�PG�V�CCNJ4`����L~���6��K�T�C:������T���q���	�m�O\�qM|(�yћ��@��̐�N��j�����Ӵ����5�1��f���a���������W��Τ�¯J����a�dW�Ж�Wsp��N� �����+����j���#�L�-,,��P LXOo��o�E>$@�@s]����'�Ḟ�7�����Lt�<K���~��z�ݽt�����r��x��ϺEm����ً��XHZ��ɐj(u�>>F�|�)TV�4&ߟ?~� z����0p�'��۠�����x�f����O�Ő*�t*L����E��k_SP��>���VG^OO�:�����6��v��B�\ �2O�^N�6��*ܮ�gH�682�a�Yd߾}�0�	��ૌғ�M�ǂ����_�45{6.Q^���˷J
+�~���'&N4��ƺ�v�f$���eGGG�C��ʖ����������ѺY8r�����솆�
�k$�l=І��[�B�G����b�q���ܖ�S�N�x��,��~hu||<�_\��:n�ʅ���~M�u/��<�r�R�������乍^�'l.T ���㾺����Rj�Sk� ��t]>6xN穙����պ��<����E��$����	����7B-���ihO;���.�j�	j,'��� �'�hN|��'X�ߌ��������u2�79�k{�p�44�����T�PV; �HB�C��@ͼ))	��!����8�n� %0�8�>7���mj��1wU-�'x�E�X�
3�g!>>���$��L���]p�"/.Ϲj3��ѩ����`�s���bl���5h�K0� ��2�D�L�ی�z����s���)9�%��ڃ��$˵p/Q�,�p��vG�H~`+����>}r@'�t��E����
K�f�M��8�&��8�Q`ٯm�NHB৥�o|-!R� �*�Ȩ�vtT%�rd�ύ}����|��X�����C�̓�P��u����g܄�Ms� ��G^�I?PSS#��	=}y팖�V�F�$&u���G��SS0�@`��lįcO���֨ݺu+ r�l�z���{@�)����:z�����6��eeeZP%Rs[��FйKr�pz�����5�$Ry��QbRSyڛ�gwA����\�S�L����o:��3Pv?���P-w����hhh��d��3۵�����[W�0�V���c��QOlA�8�K��g��FILФ���M(�'��E��*�rrr�����]#c��W�5j,�K|3`�B��ε��>J����̮��k(ml��+�
�����s�p���[��V"��ΡW�
l�b���q���v��,L-C_N,|,u�=�`�\�|<<������z��{7��UUU�:�f.]�́�V����.��R|'tx��dv� 5e>����+=�72�W��S�jfk�������i��x"�.���r��TCC��9�bRf��~��Ĵ���$���>���\��\XX�y����63;[�% �ONzz:w�jFyx�O��G��������h[p�x'��$����Ycff�j�Ę}����q�um��_���N��{vv�G�ٹ(�^��-���c�����~�|������;���ⓓ{����`TB  ��.N��n��yu�;���H�v��qt��=��*��
:����f��C"�2 �h�Li�(7���WTQYd�'7R���BCB��R�v�׌�����F�����07�g��u�0;Q ��5��V2��	t�lm�-��Bb��Ĥ��ʓ�mR��D�X�3�X6��t�u*~*9��.i$��M��,?RUU� �9Hy��+�稨�hN��@/�$��Q��\�,M��#!���yʀ��&L�~�3��?L���{����S<�bU���ʣb`s;�6����W��B�;]P�xKQ�)	���c�kv����m8�}������A�9�V��e� 5�%Tk�8���?ߑ���F{�V�q4s�z]j��!�!T��_.�����a�0�bg�ڷ�2bQĴ�������7y�sҮ����VŏY&ȱ
�U��T��pX������T�]K@ۘa�.`���`L�)�g���'1�����^s.VsO�f�_C��g343k�S91���5_C�m������u�`��Uz�HV�����z�x��+�$��x��w���?�,�#�X���ؖ�JȠtbu�~IHo��F\;s-"�ݻ���Zw30�&�t�O�K��ڼ���(ݹ��?���ջ�@:�a����nkhP�[��	�y�l����=�؛�v���kd%zG$�j����D�9���G���>_��q�
Ŏ��{�HH����;��c�	.��=Y�"�\N�8m�g��WR�A�Ӻ�0S��g@$6���w�X׋�k�#ebb�����痍����>z�}�;m���#��'�YM]�l����Y9�eHcJ����J)+7���Մ���A5f<	B6nx�n��7��ξQ'��v�~���h!нnF5���=��l��B���'�W��i�L�,��Y�ʜ��,��w�
&5]V��Igv�MT�\S�� ���˝챡���S����N1�Ǹ�wEr?�tz��2>�|��By�Wq�]J��MDp�ܪ�����~�����ѥ��dF��U���ӗ> �q���B*��ګ�β�\�;�n��޴�X��L��vG_���?�o�;����v��~���|�\���M.��<���A�����������J��ϿG���4alU�׵��v�O���906�R�&+��Vа�[��6�I2��/��^���^BBV1���n�F���e�AOI��{���:י.:Bp����6��ù���'Ũ���<kg����Ϡ����O
�Az����&{:p���L�7�ZX��rm�3��hC��A���6�7a-y_-Z��\�%&��T��J�֫��~�5�˃�k!`(��$a^}��@��lœ�<]�ݿiΞ�s����-NWgH�?�>�_8.�� �4&�o�� ��������$ r�Z�ʤ�<a�=t�hZl�0���Q4-��M%�(P��EG	�>R�	�m$mggg���f]�t�Q�IO��H�*A�#З�J���:L��P��I�T����bbu��
d�s���٭[0����d�T���Wɮ��1���־/u��a�R�Z;��rd#V-��%��*��Dg=�ͺ�U��'ƕ��D(���R� �),��W��X�&ί��w���
�����Xk"��f�4&,d�A�"r�5��9�H����ݛ<��t 6��.�n�땯���_��'I��H�jq����N�]諨�DGF���M[�����D��Iqt枮e�̲�+%1!A-���kX!ꀸ�{�	¼T����|S��Y*RS]z����M�J���6�:s!fu����ѩ��/��9v�)�]8�t���L���e���7��$��M�FV'��i)T��`���ӅJv�K�V玩�)rt�KA>��a ��r�Z;z�hZ7�Tx2�|�W%��E}#N���2���p;�&EHrZz</��J+5-��u�.:J5걱1�{��w~Z�IWA�"�ozR�W�%�ݻcRRn_�p!S�����ꪪ*taS0��Y�ȣz�/S���̧��QT5�wT��'�E��y���=���mb#%&�7��6�����d����w��s�b�Z49n<��X����(� �łW�'j��
�~��3��mȏ7�cu�Q�, �q�%���q�&r�=�d!Qg�
��&?i٪���F�,%2���#ɚt��D_���[A��PhN��Z�l$�+'�tmҩx�}C��X��@y9��h�(��;P��厪�]T������_�'Ȓ�p���?�~o���$G90;;{�y\�רycYĩ������J�+:OMn�2~��Կ/�� #��F�A��A�ɀ�y ��W9���.$��ʨĖh�!�;���f��K��0T�Y�{�O�[�{��K+��X������gF�o�}���/�Hv�a�.\w}�_G�s�`�:���1%Z�����?�dh@&T���5��H����C�������K���6;C=�*QMu^[�9}������;������x%��'��Wsg�祟>��U=oimM6j���0�t	G#`Ҏ.��z�uC�@��t7�Ws���!�./��t��bl��~8���Z�m2\LL���8\|�qd����{.I��S���tHA��_��ט&������oJ;�P?�0�d���;��B�C���6���N�8��7�b���P����t��NB���B���kM���Ҁ�!���Ǹ�����{q��Qa����e��bH���1	��Gxq�.�=9��} �ސJ���ŉx�V0Pۅo�S
[j���=깾��lC|����/�4�焄���|'�~����@(��@,~�.�����ꄸ�C9&��^ܾ�i|��I����ymW�j7{�n��]��Ŭ;1�y*�����"�]�������|��"3Ur��AV �P/��'����=�m_	C�^��
����3�h�ݐ�=s0N���)ce�$���]Lss�c�𷭭�+�3u:�t��Udee)?�	��-��{ŕ�V�T��Օ yi��<r��5n�wEh@�����a������Y�K�q>��S���@��pLW%�&��Y�H!�,�`�1��1�e+1�z������0W�����ٝ�ͤ�s�ٯ��yK���#.��(xx�`��tp�rU}�]���z��� Ө�Ǿ�N�n����C保Bd�T�v�3r� �^�<�*e�3�3��ֿ�#]�>�O$��@�srK�"��޾8X�г���yE�3Ӱ)8�C���"�GNq~������hw����Gt�C�y��}LLhߔM�E�i�A�.���H�"`� �G�_>n�ϝasY�c��s��ە�0�w���W���Y��;�[��͟����s�*�Wi���Lp���t�4(���i#ło��=
��v|���3 rj�r����"'��g�oW���p0�+Rk]����	u,�
��D諆� d@𲽃X�o��o�c��΂n�Ѻ~���4�+���N�R"�eݎDy��;�9&X��r��C�F����\�'���rRT��}���-=�z��������:�.	�|w�e^#�|�ki�^�_�+��}Ļ}�����:�0�U��n>b��%��~�'��8`�z��q�R�mieu�~k��p��ȩدGԷj�/�VE�Q�����^��z$H����~������\�)�"�Py�]0+^�	�{@)ESö����ǎ�OK=�nD9���Vf��М���X��E����l���u?��Ǣ�ƿ
���|�j�fVTTD7��\(3?$�D�K��SY�LK��H�G�OaѣqC-is]�\���%�{A�݂
񧡩1c\�.ҳ���.ں�A��߫��p�1��F.Kq|����4�^&�<j��&%0��Dı��S��Ggs�����؈/̥���_�v�����;�]�LX܄�>S(SJVgִ�Ǖ���Є�s��m6�x�Z��3ӿ|12��I�gJ�%`hl�T���AnSb�\>�� �F�\�d���K�oP�WݪŊU�Kc0�֖�Բ��zً������v(�Y+&��?��N����L۵�/��0�ݙ�����ycF��O�vz?���hn#�����>==a�m���~AÆ��Jؕ�Q�8����֦�D��R^Q1��D3�ܞ9�ৼ�L���^��g����b(��_w3��4%��MKK;O�i�V��P�s����3KK�.\��2��x�w'�X�*��V%�qb�<=:������~{[��u�+:��)n4ջ��ː�k���B�+������*R�X��\�e[[qa%0�vCKd�/eH1��c�����H	�>cl<Dΰ�
Ω�僱.w��V�;9]� ���,ME°�C�6ﮏ��'QއTU?G埐�/�Ȝ��+\��X��w2����5{����hH`'g\�E���zg��R�ʕ����������+�q����{�`���U��Ѡ���F�k��ms<ވ��a�C�o"�.�l�Aq�����,x������w�ZU��ɣD�b���Kqo�e�Fw�9�A�m.���0�N�e��*tBG��!F�2���c)�0�?�K:Q"��ã��p�8\Z.�XN�h�S�(ݍ���V󠳫��\}����d�5���i�^j0�tk��O�S�ŭ3�a���p����TK��;���|ͱ�P�2�\�̊kpW���U0�Ĳ2n]K�c/p�ى�ۣ����m��z��I���O�ѓ�4eZ{��=��f��"ܱJ��lz��(O����Zև�j]�G��v�mmB\���5>�2X�Uo�D��`5�� '���Ғ������Bw��� ���z����IA��s,������TC��o6R����ʆ+:��<��mY���2I� J���fV8Ǌc�a���}F���;��f���3Hg�]V�mw�[�3첏|��\l�t���w��߿Wo�Ud�������k��?[���Ww��o���G��!��e�ZS*�.�͚��T��	M��u��Hu!k�%F��,!z<fw�Y/��C�0N��imW�b���U��YvLI�~W����ꭣ���?Pi�	A�k(%����;F:D����nQ�;����y��w����r��3s���s���Juuu���  emNXbr�x��ߔY�&j8Z��/lmm��7�����$CI�2�A�|��h��]ώ�kr�Ôp�0�V7��v����c���Q����v�2���`����u{��_E�K��Z���-�}
�7��\>�ÿљ�s�Y4��{� ����!�6ݾ��x�m�2���H@����5�7thAE�c������!�<0�x�4r�2+���/~�|	�W���Cyטx��3���r/���$	�������`���wA�����.b���PX_��n`�!۴S�B��Y���)x��T�]�>���K��⤧����2]���f}��Ye=��Mt[����<-- ����![K!&� ��r���0,���[����W ���.h��M�F��Ѷ���Ty�"X���ҟN��-�*����������a�������sc�-�>�.
�F��[QK@�Ƞ�hŽ��c�Q,r�mu��X�}}]�cî]��8-�8��N��~���i0���L<'y��,��7��RR',����"</��^�S�U��3��uVPT4b�kE+����}��R�۾���O���D����{�AH��~��b
�d4�8�@2�p�!V'::ziQY�x=|�7+�Q�χmP���+�������}��"4cc"d����Z>k��Ge�L���N�n����r����^�z�&��#�\w=�6��a�8O�yĴBES�7U����l�}�"�!��0�W�1�����1�;����P��\��Ґ��򭍗�0�A�U=&���a����Ͱ��/�&��_���ʽy���%��a����
�>U;�d�v�{`��/-P_5uu,e����L>6_������Aae�j��r@e-����~����d5Wn��sc �b���t�b�W�
�c1'�,�ڡEЊm��43\�C�*�[�u�=� hҚ�=���qm/^�W���C��4I�Y��m���n~���<�$ro_�DB@��|I�T[r)w��ۣ������"u�P�X�ӯ�N�g��V�'0���{� ��[\\���l���:��i�E�յ���d�����7��myz��QkK-l�K�*�!����X��6.:�e9����.�G@2z�4�W:��:���ro�c�KY�QQ�u ��0����]�l�?)��r��cȴhUR��#�Ʀ����e�6�\7"�Z>����GZ}a?��o�n��[x�B'ݔ���b�[&/��q&#:J፾��/+��5j����C�?܇LUkO�*W3c?��T!h�P%�7nZ�ry�(\j�(ǣO�)�&��z��{�������s*I���AI�͒&u����Pe�i�m��&�*����<���ɘn�<�$?�
8\|lx�H�n���'2�:~��\�|W����A}��亁�Z�j5[N%�_¤�%���4�����S]dV��� �v����R���KN�W
��R�-qZ�Cݡ�h�8g[�G?ܰ�/���7/�ӑ� P(�M��-7pB�!�u�?>1!G�7�OLL<���os�����}ԁJ:�">?#��x���>᠍y?:9�3�X{!����laz�+P U��7�v�G��l�3��:�Bw��z u�V������I�� )�����T��u1��� ���2}F���4E��Q���Q���~����"ޛX���9H��6� i�<s���%�� ���s���Kh�'Қ�r��J���8|y�ݵ�Q?J��4$��3IѪ����!�6/_C���*sp�O�N�'$$<�e������uH��g�"&(�sP��WW�n����}�	Y4��
�s�0���;e��"���t1�9:��`�0|�֗㇮�Ӈ���;<N�2���m��i{�9�lP�s�Q�3(X��0b�ߵ�]V���P�tE�B~8V���[qFe�5�ѺCb�φ�O
��Z����D����дWgff��Z���;�|�O��شB.�:��=���xm���k9+ʁ3�Ѫ!�T>w�z=�����9�3�lp_�-�A�c[�Pd���79O����W�@W�f���q��0��/=��O�Ѫ[\�۩��GM<�^��F���.Q�G;�b�rY)�����ٌ�㦙I�~�3��U&����=���2��>4�
�}������|�1::j�5�%��c~s�w~~^������ܦ&]������������H��8KFv�pv�i$���MW�M͊��4�O�Rk���x��y(���&������q�����E����֦a|����I��0j�(O<\��^w�t+���l"�7�ݮ=vr�N�22(�{�"_а�?K�񥢴���P�-��0=��ď3߸���Ӈߚ ��~_�;FF���XUh����m\�ɊMA�Y����K��Ǌ�������f��i��4�$�(ʼ/�
��A�W��3����gY����nϾ�mk�'ə�H*0���@������S�?ikc�ڵ"�����Ke�c����� �hr
��߿��P�L��sz���t�{
���Hr�ʈ�T��~�#0&e\��Y��]^��;;���7��~�������_P��/�.:������A�'K-�c�d���AJ�E�Co+�7�y�&!h7�g�1�^Ն',C�u�~��_	��_ܚ��mO���]u�s��sH�����/��s���&�G/�x�՗!��'��R��eNN|O��$6��G�>�����IQ��Y�J	Sӵ����G�`	m��딓�1偭�|��g�h%�Z��)C���X����q�{`��į�.����/cO��գ���!�m�$�۷X�L_ME��HZ�Nn3������M;��(B֟��{u�+,�S�-9��b�~\b1���z����m��� .\�U�<�M�&r��M�w�m�ױ��	��: G ���]�xƘ����l/�揷l�U�]�G�>AXN���Q��Ѐ;9(b�&��-�m�htB��r3B�S�'�A���\�w�v���?0pʪ[�7�a����&TAʨ�(�F�듲F�ҽz�����
�UU!l�N����}���}�kԈ4��7���nk�t����}_7�j�;6;_��*����XX�[Z|q�f�@@�#G�$=S�>a3~��0����L�~�#K�� 	���;��6i��M:7'E�:�n�"HJv�2U�ZV�� -i͞�o��G8_�`�?���? �os)���.��m�W�ڬYka.::��g~�~�U��ǽP�xD��J�����~!������[ɟ|2�7=����ﾼ?9m�C���}�$̼�.fXv���������ս-r�J'����3rl���M��K*ey��X�#)ejR��cS��ί_�q_��7'���$��i�'�3l>Z�1��$Y�ͯ��������G�Ao���|����M_'��K�ʖ��̦����Ș�7���h������Ûc?AZCOO�K��̀ ��%a��6vvz-f�q��F��y1B���"hhF�@^W� �t���#~VH�w������oIU}ܸ�B	&6�퇢���,��Ć*I��.�L9k���Ё�� 
�_L��\�9Z��\�^0��0�3{����B��M�	53���]�v�'����{J_�����
�3$l&�d�γ�^5���;ԩ=yXه1g���.i�����W#��&ߺR�f
��=�#�����S��hS��:(�c�z����k|���p�$F[�\�8��7L��Zg$$��T%�;���!2��(m��a���iA����o�zqk:*�I3RQ�f�I�0�>䳆�zY�Ȱ��Y�C�O��>�]?= �[�3�ܐ�(rl;����~���z�n�A�n+|���`b�� � ��?M2Y�_"�7Ra3��&�dr٥a�]g��h�[znJJJ����7MO��TJm.����h�$������e��@H{��[S��\�\�8���l�̂��wl:]��Uu�__�9CJ\�}����.�9�)�f�ŏ.&&E�Z���]��]��?*�0AK��+\z\���E��a�0n��1�����X�ǖ� )7��rC��������(�fLH�'�-w�M2��
�,Ѩ�.뻬�'چ'�y��Xz±��L/>7��3�&ȷi�5����yʗ�4!����c�!4��z/7�O�V9��K�����߾�%�����2پQYI�ׂ�g+�b�lr��/�#K��v"~��*$���i%�3%�*t:�[���Y�\�݆U���ָJ�BrD�\b=N#��b|�Iz'�"�τl�I}vXfIm Qo�pL
ҡ��@BBC9Z[oC�u?��7/Ê}�~��~��v^�?��&��ς%�;�F����a���/޴-\ʇX�5��a���ӧʚ�߷��u:���ݝ�'���� 8���W�^��Mq�δ�	�NnN.0X�WOYr����d#q0q��'6��|-d.����>�U����8<L�E1�[_wFǔLjv�Js�Kܳ�w�����pn����<��V���7褓��F,������wl�sk��3��9��VT�\�u���smoQ%��W�~�;�v���ٳ}��u���hyغ�S�#��Ȑ,�8����F�[��.�jK][ډ�"��@�7��-f�ah�/%�h���斖������}�/���f�d	].�[�27Gb�8̡��I-���}�$��X���e�H'�2e�NY�m����1t����^IP�th��$[��~E��etzqw��RӿaMڸۜKJG�W��[�u����T"$����<z�V�)z�Ns@(�*�0Fr����f���s<AB��PQ|rr�t��f���+@�>��[�3)ʢ`�S�C�d��fOb������{�}}}���4ٺzo�����7�2��%�޷_�ɹd�����$��h��E��g�o�Q�/���?�X��H���u@)O�<���^m##cs��"ܶ���^�������]�-��w�8f7d$S�%J V+?��)}�vwۺ��V�,�Z�����G�~���>H�DS����زކ8H+�Y�!�r\�j�3� {�3@8�Gh�(m���m(p����Zʬ��ȩ�l�*�J?��Nac-Z/Ts�D<��s�=����0�\�۬Ө��ӯ3*��.��09�z$�\<|��0X�Ar�����\���z��t������*q����j�j8��� �D��s;a��C��S���\�����%����e�5i�5����h��ܱ���<^������E��.%�#m*��wɘ�0���p�-����f4���]m���*�HSj��k�����H��}��ZQa�v��%Q����*�k���=��d�)-��8�|xshI"c]kL�R4�0Q5��i��2�Wn�w��W0%kƦ��܂����sA���;������'�v��[���|�-�X��N#LRSAH�l� ӥ�VX�����7���Mޘ(�J�˪I<�=}:�5R���<��2�\Ğ�zU��V�<;�ڛ��4� C��uZ~�K���:4<��Ca
o� ��[Ty�6{�^�S��}�/��.*UW/�����0���Sew��~�D����/_^@z�)�Q#"#��_B�%:Q��p����_�nw���O�?.��&hr?�f����Ar?qa*0�Ї�|U���=M�"��?�E`N�����>�)�c��I\i_��V��oy���B͙['��_�T�#�G�+xM��g?�<eG*ϣy�5����e?��6���_t�݆���}�z�$�m�'���8���c�~��
}��n��#��q�z��ȅ��;{ꬭЍ/��WK�&�����(f�Pjd��ݣ��jk�l�
`'Ҝ�����J1z�K��x36r�/9k%l�ƅ	{��!5�Q���M!!a�V�Q�щR���V���1���d�E������%���Bf��$͢��K����F��5��������_�h5�,��Z]]嗕�

sp~��1�\���tИ"�n�=�Y{�!P�����&�OZ'���a�}\|� �@B���L��W��.���Ϊq�?1���c7]���LS6��,e��fMU={�L e��ڂ'��)���[p��#�hg9�h��z�0�W��ZWjL���`�����q�@���g+��V��5 �b��� �:�U� =�W�\��Od���Ba�h�ToǂD�IO�n�^�d�����{҉?b;�&O�	�3tz�uXh4����o�*9ss����� ؔ�������d��B3�T�6��-,��ѥ,��P`�+++_y��x����g�܈	[j�:>�I�}���)��������87'/��`ӭ���j Cǭy�z�EJ���2&,�"''>F�E�����}��m��R-���w��ӈA����ܕ
l����l�Fۖ�d�?�|�)C�_A�����?� v��ߢ�9Y
�����R�:���~�n۾Xl����gZ!՛��������e?Il/���i�����=
3�?}7���X�!F��b�ѥZ$4��Rk�OD=$�vи��U�}g��~����j��'���5B����V�b��h!]���򅅅2����R0�:�������F�J�nάp�y�@�7��̉���G���L];��/~�EײEu"Ve9�@C�!#'�3�E	�C�Z)A�d�����8���Mq�d�q�c&ܚ�#���a�����>�0�� |�x��4�o��a�A0`�eD������u�
�܌>.�ԉi~_o�����v�AL,	�'4��F�[���l�
Lj�X6E.�T�@h���� $
��n9��3����(���#Xy��I^(��,��������3�E��d����;6~�K�k��P&�����p�[� �J��m	�/E��NOk�n����
�c0S�i�m=�b(��!������t~ʶ.���eo�)��sj$���R�p���e}O��Q�����M?P%�ՎK����e�4lrx���N{ڀf��)����#�l���fY!���&���T$��X(��Jb���R�(F���yf��x�b?�غzZ'����F=d�=pi,}���@j^C�L})S,� ��5���bhG'<�u��Q��#��п������~R�-]ː�{�:��F��^��'C�B������ͦ�-J���y�,����&�6�D�����?�jc�΃�.�F�B�҂���^g�v��S
:��F���3Ј���"t�55�띌��<e@醆Ry廫�����f
j�Ʀҭ���-�T�{����#��WؠSjDDDeHHH꿡L���뻱�T����5f���-"w!��W�I@�J4`��O��Q=c�%D�k���WV��k�Bb�(����˃��=E�8�K
�f���
�S�q��-I*��l_����ȹ�t�![����q�~�P\_na\�Cqe
ԍ����! :�_?]M�ȭ?� ��n���?	D2w����l��,m���]JP���i]��2lC�
V�V�g���n}jr��]����"oh����Z�j�`�h"b�����f��Y��^a��i���͛7_E<�a��-�:�Կ���҅�x�u߶���-�������i۹DsWT���{Ci*���~3��U>x��" �2A�������V���7�R�.H��O�P�@�akx�F������ϼ/6¢��(�0�9�>�hx�?��ۃ��1絜t�����g>��_�ꗿ�?��!����@��i4���d|���lu��rRd�Y�uG�u�M�8À�ak���^Ӕ���_����]��M�;��p�A#PXj��xxZa#I���<�.������Ic��w��rr�i�G�v#|9�̜v*ފm5��L�*�׏�{f/�J !|����|�	��-�����>u��緉�22&���*E��%X^-����'�=�Ė�4��e����}�IIIi{����k�f>56BF����m����Af��kl����U��O���4����?�y���cIe%�\�ch��s`b���X�>����;�u�t<S��yg�TX�*e�-����1�(�Q�z�k5��l~ҲEQ�j}�,��GR��S���Rv���J�W{����J������Q�S}�S��쀈*��-[�x.%�Q �v ��;���/%s�����8�@[���:�M����"�Y��6�Mp�"^IG�V����k�n�'���t.�����%F���42P��KH<�M���`�$H�
l�����>��ҳ�H�qf�+#��Ֆ����@�:�����"���Pa> ��)�h44�\b��^qp�ZYկ��/HflV�R������`�#l���1@Q�ۜ���7c����L���9�&a��\���^�w���g��L{iQ�K��A]�E#��3ϼy��U�y�v���<=��:s�Qr�(
�6Zä�.�O�Z >V5̊������ ��}f��N�♏�"���k�)'���\��lH�R�!-ok��@t�����D�ݢ���D����eC�j,�<h
�)L���5\y)�Ho���b�\/	���Þ�e`c�
D�!J_qc��洣3�oA"c���@UZZڗ�����rI��Q��Ԛ�K���dx<CG��Ɵ����������}�b�� ����OKG�v^�7�ncgםĦ;<�GN�2���W@�z[�y�|:+[MZ���36�h��~�E�=rWE��c׶0�dS�NI7���qkrb�)~�BS���w���ޤ���0ӎi>�B��Q���0��1�;ie���2��S��Ӽ@�A�,F�Hz�ΠU���$5���gЌ�($&u�����^x���0�kNi�8�4%�05���s�/��1�����%��ߘ�9RzȖ��r��wf�dN`���A�$ � $����c����w�L�l����_�c��ǟ���ή�@麰/����z#���-:::�rYjF4�%c#f׻�dg?�B����&��J��)p ۰�:;T#�o�v5I�Z��hO܀���������'T���c[&������Is{����g���4�ǘ�7[]��EP����uj�|�E��K�}���U�3_����͠y$�Y(J&8<G�smpQ$8~��">Q�v�D�t(�g��11b�����'��G��� 1x]\�}����A�N�Y�fx8�`�Q
��������UG��tk�sh��P���L���I>zq������H�9�8#��: �b n�=��*u��ߣ��Y_2|���H�p�v ��WG� �Q �����_�i���B4�$��mfwoo[_V�#��Wu�B2�!=���S��Q��j��a�#���9\G�wYfH�����]������/�+��%��Z6Q'���S*l���I���h�V�[(�˻W��[H�H�_�ی��QkSyy9y(���"�]�Ӄ֯��ՑϞ�K�}W�&u/qQtvsg�분)�r ���F
�/@��9�P�&��L�Ǟ��`�[�s8@.۵�� y�tdJ��<e͊W4���:��-@���l����r��lM��q��]�ީ����� ~�.��b?c�յ���rJh:$	��'��y:�&"B���,"L�M�0��=��=�gl#^�(uv��XSQ�����X�s|��S[�	wo4���c��X/�*؇2Zbw��9�f�2B5���[�/E�}�8e���+���������}������E:���f���4��.��/Q[�4֭�����C�9E�����K�ab�2H#=H-⇨B�h ��	6�g��1V�V�['\@*4L]ӑ���r�7�j�\ՀT�NGj�O��&@���k����i�'?�Z���B�{��=e�|��YV�[�	П�`SF�GBqoò��i�jk/��*�����@��礤��zzzԉ�/!����j"�uo��#kO�����
������911�X\R���;{Dvи[�����2''��xa��.��EW������7�hx3%�����!x@(�r�j@���j��J��ZT]FG�Fi�t���/w�b�i~��O*�����Jw�=�hG{����Y�Ͻ�u/��u_	���"�L��ފ��oz���J����O�����:�<��{x����7�Sō�-���&
�Z�>���3d!.�\�&�5̯`���o�lS�6�E��0�PI�v/Id�D��4�cϗEId����u��sf�m�*&J�Z$�oP��k�|{NFv���'������ zn!���"vc��GK��,�s.`Lp�V��g��Mp'�hxy�ⷶ�� �яFH@�L��
3��H�=�� 7���e��dL��o-H���K�DIT�=k$h�h�L�������I�ys1J i�{��f�������8�������L�`d`iMxԗ�+-�����1���	�`ʴ8���.�T� -꯰r��Y�ܻ,4QN�_���=p"l�������z��8�E8�Z�,
�r~i���I�'�����;���ˁO��*;j�eї�^Z8���	���}�-�L�<�D����a#�f`oE�;�������GDȫ%p"���f�؛A�c��X���3����� Ӆ����	�AJ���h������"��ww߾|��9b<k���ߛ�� $\��2�5��I�T�&4�)��׸��/�ß��1�d�ќ���?3�n�fN��gU�<����_}A�*��y�3�<�	k۸�׋�첈���{�v�b��џ�Fw�"�EY[l20��t��.�Ms���N3���$���Գ���Y�/1U�1 }1�gl=	�汩�s_�EjKEF��H_�p].�k��_��/��VC��#9�G����?wbH���.G&���"[MD^_?=��p�+((hj�Ϸ.��Pr�P>��sP��@4\#�X�+(�fd`�v�@z��qfgfFh��w�&H��v����]���?sc���`���������NYi���*�J-Vx-���H�k�NF�]��E㈊�*L>u'/|ӟ����'�4Y�z��n�4ޚ$���I�����3偀�}Gʰ}.*  P��� �����+���p���|H<%Q���d��Ha5��"�s�C�F�fX�	��-ݓ�^�#*��=���m�jA{B���a���������MC�_mD��F�Ksma4$�k�Rnd���A�Ń%p�d���F�Gw�����q�Eq�?�_�Eu����hZ/F��W{��-*e׋=m33��q͛:Iz �츸�@[t)�"d�&)ݚ�=O���-�X�8���<���Z�F�MIM�0�����B��:k�l��'{��82�,�%��Ñ��Ri7���Ņ��+$��גr��ψ�/�'2>�/����VDQ�^���*b���
r�q|�6��![m� t�dhr�:��h���XKǏ ���B*��f� Δ:;<�͝�N�`
9�,�O�� ���N�?`��2zC��㊬Y�~�QȻ廙;}�?�$� .z�@,	��-��u䝆��$�w����"�i#9�Ej��888�J����8�-՟>=137w�g���
q?���1N�ߧv#www��Y�.[�V1��Bᇩ�$�o�������Y�����8]kO����P�[ʇ�Y�C\Pk�w��+�p�<�M��)��X�B�hv2M�l-m�7
�m���nnM4�9���X����^vC�v��o�VG��-�2=�:��	���K�_Ҿ$>�@*­��ÉY��ds�J{z�����5Е��v
(�f1r���?�<t;n���2Z�	���a��c�S��H��9*�8��_�v'�@���o1h+jh��� �ypL�PB���~�J~w���-2���D�s�k���>}j|wu��_�|QŌ���B��zY*w�=��S���Ժ�41x��� ��\��S򯮫��,
[2r_G؛�"P�#�m=�|�=�r �p��9Ą0�� ?:��5�'������m��cf���|�Ȟ٧���bGF��{K�
t'\���M$���23��2��H����2-4��(�9|�����|�F	`1���M���˼��~Wj[�W��k(A�f��f?[-!�a�bc�F�壸��?M��&�wO�+��\\.N�9��xT��_i�-���[��B����'8*LNZ�(� fӡı���OΞ !����
q������n�22��B��;�c��|��#��m��L�� �jj29��jjc�Ilk�3SF�F�����.QNd�\$����6<?`*l>�O&N�|͔`�+K����YH��p_�ݜ��ZddW1�M���$��~�猅��)[��y�����M�\�@1��� �: �9�O�wǓ�dCqM�A�h<nV�x� �x~����y��~e$�_�Ǔ�������ϼA��~�����]kl]�+ W9+��=���+���者��9�Q��i�,��h�w��ʾ<�����E¹&iu�������*ƛ�]ԧ�lV�rq*��KZ��ו��$��]�w�����y@ˆ]E�b��9mӬol��찺�
����A��n|jj�����F1�������)|�2��K;+��(��̄�5���O���%EhA�����s��l����;Y�+����lM��Ͷ�n�>fJ����|>ˁ|I2e����ݙ����3��?K��|߽����>[�O.o�k׎"�W�B��F'���0<9�*��)}����3�x�����-��i�'f�&1�sχFM[��������:��A���n��qx�)}�K�{�6���,�KE>����bps�kG�I���weҾy�?���($D���*�Xb����Y�?��Юc� �>�
�0D��GtJ.V���o��輷`��-�gA
�,�\7��ۀ2p�Q-���r�gd�����X�	��	RDs�j9����VY�%�9be����U<�}e}IrE���d��Ɛ�>�h*����:�/vB�z�����#�N�o���[Pr���OѳI��8RS�g����~{����A���G��G*/q��ُ�%�V ��=>�$w��8���_���\2�cO��G�:�q�Z��;�r�8�C+�����T^@��	�s�l�]I,����-R����_}���ܛ0�=9J��[��y��w)�N�f��L���3�M�=��F�r��d���8}����o+��Կ�i�M�Hb��M�c{���c .p������YYY��q~(�UZ�+��u��09<�*����϶�daS���CBB��������C�)�����.�����e���dQ^�_�����"  �g��m\D+��_�=���f��X���a��=��
/�,$����5��5��^�����^���ش�z�"����C	���2�Zj���7%�S�њ5x�BQ�vW,~Z쐍F)Y�՘���t��S!��d�{����]���e\Y�����D�B_n�����۠���+�]���U7�l�?U��%�{G12a7�������R�V��ϑ`���L�f�:�u1��&��o�94n3 ��FB�ѱC�P;�x�NSRRj�)��᧓fm���\gĳ�C��;�;99��{�J�ݞ��ߤ7���3[m�t�ď�?M��ШI8�V���uYY98�s����w�e��<��h��[�$�T�⭳��]yxxEz�/�ӧO�63s)c�R22(�-<T�{��^�Ō-#�ft-[�T�*L��ӂ��>環%�0�=�!�~]�~g�c�f���i�ܣbo��Hؕ���aiۛ��K�F~ k����G4ʲY-K�Rgvz�6�8��yN��	�+)us�͝�ö[�Ei�A_��>�Дh�q�1��r��[�S?wƩ(�.t�� �����]�^�8�'e���Č"j�I�uWLrD|�PÏ�D���$ �&8��B���৯~����oVI�K�j&ͱB��Ds7)�R� ~̸��ߟ"B¨��S�	�mXcB{{���$ߙ����<Z�t�1|�A���#��|,c�X�@9����od׆�H!x�r�.o���8W�[��J�	�> ��Ru�P+ޔE��R����u���m�`��h"B��-��R��� �%%k�D���&�Q�!j�3�����v�T���Pճ��l�$Ѽ�ZHL�h������.郾:�r.?��.�G��tw6��t"2_�B	��ow���ۜ�W~=�,�h��+���M�H������ĥ����`я�����p���i"���o�mo=���-�-�p�_�D�5j6�D5��f�})�,�} �Z��ߪԃ8�ی���2z�Ɵ����,Z@Ԫ���ҡ��Cn�tTb����8�G�H4~~~�@��.ќ�����8ۭ��Q�ۂhDdd�㒘 Es�aЎY���in��H��' ����4�P'0�!��Ws9��U�^q"A�����a�Â���"�B�U)Pg&@��D�W/|�(OX�Z@�ά�U&M�@Q�dR9o���K�8$eo��� �}��YK'���aP��U}�b�'y����L6������;!�v1�ݠC��t�^�R^����չ�JQi�g�:��=�'}�п��Pn�nB⧷����'���P����M��ʝ��Fy"g�De�9t��>�,� �I?��_��-���c�h�{�����-ܡ9A�kA�����l�E�U���Av�v(����� kp�/3?�A�`iaOѓ�����"�ǄK�d�"��&H���3��eϯ�+�U.�>�"�B�ܵ�t�J�.W�����C�b�WO���I�'�%��E;*Q2�?4�>�D눋�>�F���ES�G���H��*Ƀ�F���4�~&�(�.���;]�Hmǟ
�����,@�Ӹ>�Y�৻(9�.==�s��7�-%꽮%"�p"��ny��쏉��%��o�=�X�@�d�� �t�7ՠ�&�E�Tid���x��N�;dS�|;D)��8��9nf_%�'���7<�!:�/ �fp���2�0_�B/$�W�Y���مσz<�FK�'�B5�`�1�~�"Q �)�$a�8��Z��g��':%�0�X��;���+(H�`��F}�X����롗�����!z.<����Fp�,��w����jk��joA��za$6�^O��g�^�����G����ԦHhC�t�Q�'Y#���(.Zچ
>�/5Gﴣ��m�O��-6�q��W�E%�S�!�.s��Z(���N��?m��B�w��ڋ��%�j���/y%y��BTgH��ڶv���K�_�r�I����l5%�l��U��s���Jn��z�������6������{���#�ÿ�A>=C(,,TQSQʇ?��2�5�0�<Xt��^*�y�6�'�jE{��H������Y���\��T<�-�,c��zG�p����<�,D�x���ӎ��gu�R.���ٺ�$a����+��,�[�>H�,��<ӹ�`+�o�8�`(�	=Z�������4w�X��Z���B�ʨ��9u*���R�τ��4��<��5]KQ\������<�rQ����)؛������?�רp3.�Ӿk��=j6��t��j]U財��;�%l�u�t�w)�M�i��RS4/���$ɟ���X̶�Ø�J�$��O_�/�dA������T^�	���|�+\�����c9Bv?y�9��,�;�}�2-z���YxZ666 څ��~���r~m�ߒ��@��1�,S�#"�Y67~d�Ж���'�ߧ�:���0�L�d\�����iӖ�Z�ӹvtq����2�E������-��Ԥ�h�|Z �a'�3����Y�#+����*ֆg���B�G���*ݼ�,_Ms���u���n�5w�w}�tm|�����_D�kz�4\4=����JZ���`�_���C��$����$�P싃���K�����ފ�W��R�_#��z��nymln҉�REJ�Y[0cj_А���)���d0( 9������n%:H�o�~���3�>��x�륟���F3-��Ĵh�t�����/DXhI�29���l׾�cd &<�̱�3����P��W�Yﷰ�Ÿ��j�myu�Yr��Z\.��ĺ�Z~Uf%��D�T�����]o�����T�#}�����vH�|	���:u=��H��&�q��*���M�1�'tst���['�"<����я����x�]����qo���m4��`~��Zy����L�;�>����%�`�IPj�9n,N�ml��D:<�c��,��ڨ�>6�լ����y� *g� �,NQ�/���*Q���@m��R�N�M�8;J���m>��0}�W�3���!2nn������XT�F����sE���v0b�p�R�>���Κ�x(}�X���7�w��2��u��;��A鲰z;,F��F����j> n����%���o���}��N^��F��P�5��<]~{VG���kjF@i�1�ٍ?�bK��2���/*���A���$��@��	��Ѥ2J�?��#+޻����B�#s����JF{�<[�����]Z�p��qR�p�Y�p�3�dL'�G���^�m���7G��T2d*D8�"�~H���X��Mlֳ����_O��|�]s�ͨ]��V4������	�+�*Yn�!�q��`s�ѯ���h��ӭާTR��s*��>K	�k����p{y��?]��؟����|�a�/�@�uvJh�hv����p��J�ptZ��537?Fbǭ�q�bR�A����y�oT�ޙ &1�}�`?��M��W'��G:�ͬ��Ȉ6;��p#,"H��:{��O����Q-���<��!����8�8��^�ϻ��\��1�����<���V24V�bW�=^@���/9u���_	
�15:D^�,I�q�V0����ꨨ���AQ)I	�����T���DABZ�[@D$��n��x������t�q������8����,���VՓ�%>?#j���f�wW���gz�?���ܒ�Q�%)S����I4p���g���Y�8)���z��M�5�*��[1����t��ӕ<�qG����ɡ��Ɔ�����<ڛ7w#�Eԕ��A���B�8����N(�*��z����~��R�Yn6H����:��Ɗ�b�'�	fo@`���3�C�X�'ƀ�d�r�c��09{
���m�Ņ���g�L"5���4��F��\J������LcH�RD��<Jz��Y���+���a�Q�>Ɍ�s�v .��]F2�䔥���=�9�MLđn��[�W�Y��u�/IZ��7����ܝ)�$���g����V�q�C�w^�Ȕ����`ëB����&��)n�3A[�;a%qڈRΆ�����_R�3��ӏii}dc"�Ԓ����ev�bC��@�)(Ȗ���$���P<����M���0k�j_K(w���2�8�G O;�O��Ut8��U�|-b(���������]_��~s�����dm� �u�3�);���`�n��~����`����##GMMa����&�fP6ٴ�z���4>�C�6��o�q��Ȼ񒯗q,�@��Ri�q��"�s'�����l0d!��!沅��*;�T�ę�t�t��Zf��[p�3���P������b�xxw�%��7������e��@g�|=c府�@?�N�������}��*;�v*-5��Y�o�.�#Ra)���q�����у~mzb��|�8T�{����#��:)	��6{i�ƀ7� �#���(Bʱ[Uuik�3%ẍ́���c�)�q?��p�0�c-�a���!�3����g��k�P8C�B���eC��-���RE�58�����q��ʓ��c���'��(
>�̝A\"���@.��^�4bm͔6��nԎ-<��n�&�䟺��A�"�G/���.ICq=)ᙢЧT�M\;}E��x��+ؠ&L�|}u>�n���#���v<V*D�N	6_��?�i	K���"�1����5���J���'K~T]!�׾���[}�ر~yz>���8 ��8a��V+M���;Wơ�`�U*)�ZJ@v9�K���E/��(F����q��߷"[��/k�̲U<��k|`��س58ʕ���+o��>��\�@G�$��f�;^ցR���_r�}W�*�Q�K%��v�Fww�}<<?_X�h����.���T�I��3s�(Kt|dm��a=u�Q���x������L|����"�k3�&b���U�F󡷣l��î�2������",���3��ln^����K�/�Φ�,C
�`?8kwՉ����~�g�̽�Q"�^��%<&�d��u3-�L�h*���<��U��o�@���i�r�%���:� �^�����4���9�f5!�L�|Q��l�-�O�Zr�y]{+s�ߠ5��"Lj��a=I��<<O��/��T�� ���D"�65��JK;��?&$�I��y�R1n��������J쩣z�G����m1��r�I$0L����Y���̺�=���+��d$�A |у���-��*""�l?��`[��X0d��j?(iw^[yn'P����)u�_v��UX��u�����6O	�5�]�����������	��Esu����^q�2�'3O��+A~�*lGԳh�9%���4�?��R�$����FJ�#�a�>ߔ�U��L
��#/*�~�pn�3I|,,�2�--�G��9_�ES���ݷ)j��Ds���gTÍ�[��v��x��:���T�@�k6R�Xϣ�Q��%&����]�hʲ7�(�!N!���N�z��=�������x:!����v�Q��C֝m�<���|Th��l�wkw����;����n��G SA�]��}^�.Ш����-L�����A�0��!�ى��S�z�oEruT��;g��װ)�?��)f9Y}��e�C�)A��qbbb�ϵ7�*�N�Q�����������$�ת��k�H%]�F�j��&/Skk�7����X��PX��l�0(Ƹ��^���^�W��p�i)�ܢǖ˭;�2�&�vߘ2�K���9~�8h���JF؍�>N`gWV��['���6M p.ۨ�
�ZT�$l���q�멉dm�[�!5��s�vME��M���b��ɡ[�Tp������X�Wҹ,���,�i�;3���T�C����e�G�=���8~���HL�hA~~�H�6���_��Se���v;0^;r1SD�o�����f���K�n������NX��!,��UN��O�^{k��>�uT'��c��y��r�^d��w��;f/"�B�f�l)*�g��΂��[~�z��[_��Q�,F]��PԷ������5'=��e�N�M���y7�j�����p$zq��R�,�߲�iXG���	� ���/�ҡ�"�H��?(����Mt��*��/_:��߯U����A.�����Ee�g_a777	yyq'��5b���(���J��?V^r�u&���[7��m��o���Ӡ���`�{���~;�w��
S�r��ul�S�s����7+�÷�a�xt�t�n�(5��f�vx��.�{; ���*ϣ=G�}�~�#���&1-o�����o����9��x7���鷯e�p�_LceKQ��lw(�x/�Y�oߖ���`��1����5�z8�-6�Mߋ�$
��Xd�P��9u��hck8e-��n���ь��K#�w���G�ʧo�'h��{��%%�t�����Q`���*E���F�
f�Hrr@U�G�;��� _�b��֖�@+b�����p�>8Vi�+%%5���r�%��ʦmV��5e-�a�#a�p�lX/	%�ZT�������ie8m���ۼ5l��ƅ�d�[������o��	�ʘ��-���BTz�0���M_��f����if"]���h$p���oK]7y��*^D��ś�xE�E��x0���:����5��O�:"6>��6����߉,!	�n�D���`?6v�6�m,P�����Q^�'KS�����ЇJ���l���������[X��b�~�Z��E�D���y�����B]��m��9��/X�B��[���l����H���̢�
V�n{��R�R��̒j�1aI*1�<�d���ckw� �I�j�c"^�/�k����_JJ�ux���~�҈If��O���J�A� &�O9�<J2&�`�i�ܸ���-ѣ��U}r�w����Ty��<m��y-���]�gP&@6�>P'��劎�x2�^���C2���/��6M�ڏ��"��Ԁ�:f�%��p'�Z�@�Q�>#�u��#�Q����~!�i_��i�:C��E��51t3�2�o�/j�f�lx'�e�N�Y˒�}����i{���CSS�	K�|(O�3�w��*�
y�N��OM��k�~���z��a�ٓdJ+@_�0�ى =T�Z����tGd���ng#�LrVgA�����Wl��B�T�]�^;;s@]�=Q~�X~r��rX��I�zM��-��� (�uԄn�z�a����ù�MW�p��e'
w���ҽ)}LG'@���.�
 �2��\�=;h���)�U���?�z��"����i-)n<�=V5�%�a���ܐ?�'q{U>bVvh�H{�k���"�;�����W3���B"��t~��G���slg��{P��N�#  ���i�KLr#��䠤����S�۞�����P"�KbNNN`�+=I܎4���Ӿx���2�U9(��QPP�Q����`��R�5��i��\(yU��a����ߋ�w�6�����B���\������}~.��e�p�-�58x"&[1R�W��RPI���Ly�v�!2�nj�}�l�5F�07=J#T�\.Uכ��R��*���%=$���sM���iO8s>�Ѵ��������S#���F�6w���{��q�6(��@�X���k4MMM�*��ܖ����L

��"�����&�~>�
�1n�W�-s?2&%�͙�":b��_�r�L?�I}�b�>���~Q�3�v``���F�E��t&Y8��1^��	��D�!���g+2×�U�n]]M��j�A%X<�v��^{xEw��&>��5=��1��BLd��Y�O�[��@I��ӈ �C���fI��?~�n3��_5`��M����d�^#���vF$����!'V�[���쌸Zz���X&&qKw,CTJJ�e��T�===\j�Z�8-�B�DD����p5"����;	_�@�z�0z�~�`�A��)[X��?��$����^�bD��QѦ��X�\��J�TQ2[e��F滗�G�ܳ}Z����g�i6r{c;���\UG^�L�0:��IT��l��o� ���}�2������>S+�.ʲwE�$�!\@0o0����6/�v���)�'�c6�O�z��17��餅��L�ފm�%d����CEš�{��h�*��f����1]v"g��K��j�$r���/��e��"
z]6��&i��JCi}A�T�Z� �u�D�ah�}���|G1������%�vK�iߠr����cF��00r�8���M�Y�?_'*#�2_K�jG���S��&��q��[�DC�m6�U1��/�����JYo��w<���3� ��������J����u�v�C6�.�(k�6f�"����|�C�!g���ǰ��O8��W���3�qc$a�Q�<q�����0�N#�o�㙮��|6Q�}�k�b���f��Q�ר%ϻ�:�>�j(4`�[Xx=+>u�WH��d-Ȗ����K��������o��6P�?��PUR��:Hs?_�U��*�����=}p���u?$��e5�^C��~ ]�^D3�nDCt�ӱ�H�@���zY�J�o��0�����}���I�!�Ϭ�q�Zܦ
T�)���&5;֤�+������z�Nr����G擔�
�(=$l����7���VWQ!����ٲ)8��M����a\5�AUfV�co&�.-P��lQ�h�������X��w�,���������*�E���j-��7�V
iZZ����rY����6���ݻ��xߙϡF��E\x�Ul��D�`*�I���SrV���YVb��T�G=d���%��:��xÖ�F$�0���1mZ�u�v�8S�	�-[��c���ԝ�\��SЍ���U���J�X��|�DG��bS�k�u����P�\dǬ޳t}@Vg=f�7�Q�7�Ф���q�T���tzAȵ��g�Jh.�)Q��y?�"*ؓ?����n)�L��%%{���3�뵟?����Xm3˔��Q��C�1�f��N��o'�iboik�%����'�an>9s����n稈\��w<Y"���F��	!��l.��Wg�C(�򜒅ٶuK�:Jbh'�X�3�ޅ�$�+?Ϳ+64�͜8�G+U����x���i������Y7��EP*s9եz��M���l쪚n�\�o%��=�@Oy���Ҧ��EC'C�����RQ��xLRL�e�ӋL�!s0yD��*�\�\���-Ӷr�`�����u�aH���,ӧ��^U[��GUU#�lB��=|M6"U/��j��'�H~E���t�����[Io����� ��3e+(*zѽ}�����j���OUuu{Љ_g��{ނ'~�sIS��J�L������DfXEQ&v�-mA7Q�Y7�@Lگ���}��ݟ��'�e*�m"�� ��o�̊
���^G����_����7�����_T#и���k���kQ(��i��w�z:��$����]���hq�j�j~�C�(^N�!�7Í��vx�q`!��/��T��[%�_?T�����rP��r��q�E�l)`�ƍ�5)),���ЗA�)�o֫w�RRV��!w�r�NX�C9VP[AA���jltt4��oB�T^��2;�Ah��?����}��I�N�]#(KS�����X�/C�z�źd�e��P)��#�]��{V�_�`nƣ��u↤�ݙ�����u9���N^�wihZ}�����NӹreP��k�A�BE2�{e9��DkfB�7=�/�Ӿ
j(e�|/���l�v���2ő��KT8q���gS]kX�>3�����g�X9L#�/+��C_�\e�5��!��EH9WNUH�ω[AZ:���[�nu5���'�7t�%�_�]]]D�Բ�Y�J�.y������ T���XAg�����ݜW�U�i�coG�H67!_��v»?J�Q���hM�e~I������{�˂"��>�~�=g�H��j��Fas����1`a��,N�
T�7�P!	}3��]���b&1�Y���sם���]�Ɏ����8�����JCNIzr��ȕ��j_9Wf����������x��8#�C��tԮ�d��ǰo��Ǚ���2��$4�����
k�j�Ԣ���Y8%QD��I!<###s�e{.�[.��ӡ/gUQS����}y�A&дӺeo7����:1�5<2�����I���O�Jw
��3�[�Z�,M�)��=6ֶ]V!C���+��?��Ӟ[J�n�G>�gS�=6e�^w�=��͑��Gi!C�6�s�G��W4�6�J3��*�tF���d-F&}�����;%�U�J}�3XTiS��a@8y5V3<�cH�H��Uy����ƽz��j]#-���6�u2�FƂB���ק�j��چ9��d��jj�X���ӟ)~r����T�xO����˫��S���^`��M����h��r9g=?a����b����e���cP[㽮��~��$|���1��Hv�%LO?��}��A0T�Y��ьs�5�*y#�'�,����$�`��#�(}���gSV�z�ޙ��Y�n�H����on��7b�Tj��}��S���dy�t��9�g��`?m
�+�+�@u�S20��˩�Iސ�jaYޣZ�|�})ǃd}�B^gD����j��}4 č���1
�/Jq�;���o�^,��ri�'�
 b7�	�I���{�Y\,�W�~��=sSS0�wqM`0�-�+=vu��]0d<�<-Z>�wQ��.9�����y�=^��vC�0�zp�/�F�iφ>�V&s5���`m��V#��Qj��A����3��M�g��M8��_�Ṡ�9�PO���~��-�Ƹp1ʉ��ҍ$٧ �z�ۼA����7 ]]֨�i�?����SW���r=�Gn����<�d\�ڊ�1=;��c��r"������=V.lffFOO����u����yͤ	�u@�v�����R�Ƿo��9��x�i�\;:&5uFݙ��oo���! ���Gy�x(��Aj�`\r�g�bK�R�X%;��B�����=zgd��W��I� ����If�^��&����H�fw�xs��d�s�>8�����HOe>�^:)%!����0���l���IC�B�Þ�u�94*ʫɣ�ӌG�k�Z��i ,2"�o��&e���j�sw���ui�SM�9��T�^Yw8����F���n�V�xJw�\�#ia�!��֪**y�����c��GG����P�����{����k����{8'�`�I\RXXh�VO��K
Y���ZzZZ99���~L\��S�� Uhiie��=:��?Cy�~�4�Ӣ"Y�m��a=W�w�˥D%�Õt���3k�T|����_Y���ϊ��|����N��0���N�Ź>y��#��6��@L�f�s$!f��ݵ���/��U�s6gk�*Xs��i6��HyN�/�V�*?���|��J���s$o^�:�)�&б��kE������:y�]{��~��'=���\�Q|=��P*=�(ET�h9��z��/_A-��k�(Ű���MU��� +��srϮH�'�+Ԓ�'�|��w�����"���B��,����]IM-n`pp��i��p:����;��uuĎ|�a0�w;�'�@����V��#Ot����N~�:�co1�T ��v�y��6o#	��2�����Yh�>�HƤڸ��g��~ k�߭8���օ�h�y=ޥd襃��8q��@���*���)�gDuM�gǵu++4�GZ�f;�hhM�B]TX+����;�d\
�dʹk�6���nojv�R�v�O�S�?�3��QT�����h0''�|�dUUU�|���$A���ԁ(VTV^�;tu�iG޻y���F]\<HK[{@��6���+��;i0Ln��}�߆.��uv*�����~�
}-;;�j~~>p�/{��f�ߺ����\�بkee养
�[.�<ј=q�m���������/G�w%⭹�P��M�5Q�/l�X��#�J/�v���,=9R��ib��!�ŏ0�0�U��JY"�ԯW1y�d�>��r���~�A�}}� KQ����Y�'�Qf�*� ��`�U�LN{�i,TN�IkUH�2�����vzb�	&�D�ț�$'k囿u���M*��P�$�@�a-o�曌ʯ�:�̣�W�^�� 5���t�ӌsxuU������`+�����������ϕi�����џ>-;�_�U��"�/=0�]��(��HK6N�d��o��;�)AK�<��C?$�����J?���x��7�Y�9���`�7�2���k��T��:!���p!Q	I�U�h����~r��=ǵp�GJ���%��C��%TE�5�/S�=�|Z��e�s;Ҧ�Hr��̇-=�#�; ��T�=St;�Z5�w6���M�}ֻb/	p�=��1���FryA�eGr�b%�57`�������mq�����^�����h���I#ř�e�Z��J��YT���h�ݛ7�P܏�n���͚y��B����z	c��=r�z��	���������<a��'�;��?os�-Ey	��K>�o�L�K���K����}j����s����}jR�#��ӕ������7{��0!�|Y�����:,��8���!��0���$�)��'�2+7�V^��O�n��%If��� 3���,0j0TtlBƅ�c:ӷ}��?J�$��%���je����Plll(� ��:��.����:��������kЦ�u�U�k���-��ۓ�����C
 �Z��"ľn�O�s�~�^�2�pӼ
�O�L�ی�Ì�"����F�1�m9��洳�j��&�)��o����[3���D�[�gՒ�i��9|+�k�%�@l�OcM�j^۔n;����3 L��k��F"?U� �ί�@w���Zyv�L�蝖x��2�g`p��:�~(q@M=ë�Ǆ]��*�܅ׄ$S޾B��yC��o�`�)���`��Kr�ժ'��_�U"�ȅ�J{��;�����@��/%� "��X����߅~���1���C�hħ�{Tz��9p�ӳ��ԫ��v�E2�����^����O�E�T�1�g:�8P	:QQ��՝$�����χ���ᆒ휮�#����M|��4;�P��ql��� Jߊ�1����ŴK���Z��W�0�5�Q�A��U�YS��H/�(�?p,��8��;�c�95�u���4���0t����W��E3��Vc�1�Vw$�k>��6%�m�u�t�*@�h;�I襖ʮ�v��XdC�Y�� YlQRV7�W�Cw5u;9-�'�@u������+]F���T�]���.�g�/�9`{�][^.E�C'�֟n�`���eJ(x�5��my�K=��4�T���	G�k��Fi�QtX���nLttօ�7�q���s��ɼ�f��G�D�ꂅ��"��6~u/�忲�u~�|��������� ��'�5���K�F
�����F��S��)��5Yf�0�P�ȦQ[K�<���h��a��3���~@7�)hI�
j�DMq�����	�K#�(���^֖���R��{���I�Y���}K V��+7\��:cMe-��(�����p�N��Y~׈�d���$�E�a�*z0��SnFT���@¯܍J2��K-�O� Y,E�k�x���x&aK0���׃4Z|, �F���x#/��y�_.cʣ�:yc���zT.Y�����ʧ��+W�{��g?�Y�6�p����޺�%�X<]A察��gT�Q9���3�.��W=�6lI�<o��`�[qc����:��f�K\P�����#�S���ėYl�gF ��	nR��M���ɷ�m5Z�r�o��r�Ef�@�6�ֽ���Z{m��2r{�WV����ڊ��| "��o��e�K4#���6�V�˝�c�r����B&ԃ���vP�����@)�h�#���n�r� �p/��9��w����O.���Ύ�M��#/��r�d#�-����ΡB�L�}���D4� ����R ds�އ>�7Rz��03B���Z��U����3Sl���1�$ŊD<zhp{p&���\2���[�v�G*]�uϔZO��*}�Y�8NJ9H���ў��y
ľ�����{GE��S��k�~eL�̈���0�L��i�(��.�V�I��0���h���6� 	�����.V�⵭YܼR��=^�8`f�z;���\��N[���,��p�Ü����B�]�����2D�S_�E�?�6P/<npM��6/��a���zU0D`b�'vͦ`�Ѭ�3|~��U��T�������KM��C0��b��ݟ Ȁ�iU�+=�,l(�%�w�����d�Ms�rtl�4�Ga;i���#�R'�4yǉ��j�����ju@M~���H�֬��`�U�z�h�P��W#V��Wr����}�~"|��yA�-EŮj��S��oj����9�����i��M6d~K�6�g+��>}X��Ț�J�o�zw[���p�ЦHBP���68M�:�������dc0�뉳���;�7�f
���y�_3�6Z���;�xA�$�?�"W9�HB��廇��Zk��"�� �r"߅����AAK�vjQ:����?���/v�IJ�Q�����j���R��辕Pb�J�?X	�J�&&���k��q�6�3s��l���/�i�+«�.�{�x��b:��=���y�)[�J��n�%�@���Z��R�w�Ǯ7�7L_��I�+�9m*f��7nh�+Ι���d�Q��l��G�Fg./pE�����l?^f��$���M2���F��Gb�rIS�T��Z���� @y�{��mݐg^�h6���M�=�`����yI�u�h��n�4�l9��h�����V��x��ba��Z��:�V�f_�����c��p{�y�Z>�Z/���Uj�>�Q+=v?[�V}r\�@���"
�Ҵs?տ[$�,�	c��~�+��ٱ�|y�WD	������`����<��:)��f����?Y�>3�����S��9asuƄ�!j�s����`��m[�>$���ю��u/JV n|��p6?���j��0Q�8f_ߞT���2l��.�7�@9d�V\�>��g	�9! �-x�eo�Ւ��P��v�Ϥ�L��cu�����hH��x��7��J�Z�/�_�/��v��Kth�{�%�f�<�H8�4�zgů�H���T�3�J����I/7+@ 5� �b�t���y��4�p���R�pU�#����10xAt�pI��Ҧ� iB���F�x�$�n����H����&4��������Dg����E�f�l
.�:}��\yۖ0�F�e�>2�J_*5/FQ�@i�&�QX�[�沩��'�}5��U�I���![Gu{��������&��l�������V!�qu]c��A�3�\����LM�s��|�~毚��;װJ��LtT�����^ UQ
��Kv-N�kX�\����f�� CC���U�ݧ��=���tQ'IMr�P�;$��oE��!7��#�h4�kP!]�R�/��� �b�k���D	i�6^����9	u�r�ʜq2DLpz?�~% k���,��j�]�����utc�	.�x�[g�v�4z��w�ˬQ�t���5�t�$(FAk�׼����8�7���t���̘b魎�� ��,Op���IdmDtoO�9�����O�FJ��[��<I�T蜗�.b����5�S�Z3�C�C�>Zj$���H �Ԣ9��E�����O�J�K���ԭ�b9��=,-Y!R�v�V�*��yb�3#m��Pr~���E$�������
�ʗ0,Px�` ��q�S4���W����T���;;w��4Ζ�6)�vt��U�]"�W�S�U}���S8��t�K���GK���>! �?w�9��k�����*��7�k?T����kIv�NH��x���*i4���2�J��I���|4R�����SJ��k���v��nt�U][�g�07e��Z�U��^�x�J*2�+#֯;A�)&g֕��{$�@0���ô�Ù����{%
�hg��)�J��$!ܸ�V�n���NחKͳ,;7��Re��?u\6: �3���j.,��
����A��X�7)��#��g ��;v�p�3_&3n�`s��1�,�nn�D�K��|,��8X ��|r�8FY��aj���Hq�)�$ĺWmڳ�B��6�*�=�	؀�>�������9$7�X`.`1�5�Ux�Ԕ��M���o�:�}�2� v�R/T�r����۸g��h H+���zV������	���uk��F�^(����Y� �N4�?���=@<��l*�ɧq���4z��F,lu�&�������i�]� ��C&�F�pT]���W4s�zZ��׸��q��N�v�lú���F���ʅ�W<���<D족f��[t�҈z��1��W�����%�7�S^�]���y=Y�և�ZsX��gl�K�7�-�{��Lt�gZ5�E 򳍍����h��Ϡ-��L�:f��s"��_�<����Ll�����8�ׅ>=0�5��"U�r�@�7^���aC��(t�K*y�Q�x��.��N �����E���j�@j�N��5�)�M&�@J�M����<3m���~������bbh�q��dQl��J��厡8���%�)�<�I<HՏ��������$Y8ϱg��r-�/�(&�
��~�L��gS�O
*$�+���eAd�����gc�zݺeP5�����)G$!���~��M.5��&G�I�5��{n���{>�\E�G!���U�U
�&�`�AR��-JOd�a�jh�$T����ב��厙f��"�+M�a��.����� ��WK�/�&�3�?�l˴�KQ@��]�tzMI� Cg kX���$�8.g�؜�R���-����D)=%��H*�QQQ��-� ���*YKO�[E�N\߹ůF6b�A�7��豹<���E\���t�(���y�Y�)U��j4,�)Ԯ�݂'ʰf��ĐVy��a������GO1�SC�!F��"P�������~��î�����'�k�5���_8���V"�/��:��9	���7T+5�a�.��5�W�z���e�� X���:�K%S*��$7���"aAab�����<�%+��"���s���*���m�G�iw"?�,<Pj��~�W#X��g+�Hym�"��;�&;jl��F�(�\�ҥVw���
�乻�z���8�������dҺ��TW�y��I������=�7��-pA�a�� y|���
'���=�<�=��Ap��$?���������e�!N▜ץG��wb�T�z��35���	��c.s��^>�@3��avG�(_�:�(�J����H�ǋ"��3t����S䃀�����K��} �
̠�}?ac7j��Pw��/�t��1�u�Z�x�&�8�0	ƗF�/%������M��J�U��jñ�Q`��M����l���黷�vԬ��'�>;~g�h�˛:~?me|�˴���̞�لN������&��{����K-�p������q��E`�Mє�ab/ ���0k&���.���s�	�9ТK�ȍ�� �N��v�nQ(ȞB����S1꿒�yAH�/���N�!�C�U��E˃�`�>�Ai`ńDx���<J�/�ږ�^1�f�<)i�l��`���J�o3�T��j*�0�S�z����hv��)G>U�/OK�C��$4�ǂT����9e;|G�sY�b�MY�N��"�G�eY��@�#?�����3�╲�鉍��p>@;�>�?e�y�A(� 6�hr����)9z܌�V����c9�����R;W����i���p�@C����I4�b-;cW��M>_�y@c�g�H�x�b�4oP��#ߎ�����{��Cf����Փ��?»`܎M"-G@���kT�ƌ�"��� 6���K"��ι�����lKQ�$M��������������L�Z�
g�c��1bC�Xڈ�ΘB�:S-��"�}���y� X@K����y$����SX��@�ēu�A�X�	Z�B��)�\���?��l��S�������3e_����Ú_mx����H)]d�T.s��D4B��ɗc9��< 6)��?�,]�ZP��l�
�y߸�m����A�� ̀��Gr0�a5���#[���4�?����qH��I��L�-#��Z%�a2�w\�%��*ۊ_{�~�TQ�h���pDa{ �H�U�R L� ������꿲�jS�uxq�:�ul�3n\ž����Ti�
^�d�4���&��밼'e?齸lK��2��CL�׭��dڦp� )IɁ��������Z3PK����D�5��Ŧ{ip��7��S|Vd�0 ���'EPa�<�e��b�����A�0�Q�Z�������҇�r�`���������N�vf�6U!2��7Y����DJ[?�ww�2� �{#��)K׼V�&�o�0�S��D�g�Z�nc֩4�b����~N���_�J�~����ߔ��V���dZ�g���x��Af�Ў�;Ku�j���"���ګ�2��̳6g�Y4���S�P��s�0��Ŕ������WLH�`Jnʁè����#棯�`C�W�6Z�Εgп
����1�sЗ�%��In�y[�^ǹU��O��P���FJO�R�[��O~�U���p�A���P����#F�:�`��+5O��f��g�᧑I�i��� �cIu��ۢ��W�/�ð�c�.[]6b����>، r���*�l�S	�]�
�4�;����]S]��G�{�b�ޗk�O�	��>'`��+�L�T�d�
,&�&����`�q%����I�`�eY��V�������Sq8��t�n��wu�J�B6���Ө|+	:+'�}��o9C/�{�U��cA �]2e�!���d�宝�_���lIU)��ܓn�4�>��/k%yr�,�I ԍ]U�J��.OJ��O����7�2;$�����,�R���\c���{Ū�~�MH �+y^)���h��8�6.}�'�ݼ�,�����f�i�����#��G����;�Hʦ�6����B��w�{8�q�Z+�(W�ڷ,�ð}Gas��t���(��
6D+o�㳢Ξ�-5p��o	�#� mܔX�.z�6Gh}Ʃ?���F�߽ٶ_�aن��O)�W���%�̈́���M�H�.I�'Oa��ɭ���߃)�q�֣�8�ttϧ_ ��R�3��C ���+b���zj���u/�A@���џ�y���ҡ�u��>�,!��X�b0��>j�q>�����';�q��{� �a�
L���W����D+ye��J�^�%�&dԲ����pE4R�#�l��L^�FE��	C��vg��O	����o�(���P������p������ �N�S���w�랇�)B����{�,����}[�4Ö>��y�]>��1�����=��K۟qd�Y2��R���i&㤅!���yǻj�ŏ5Mp͆�D��Ͽu�|���sL�Lβ*-����΃l����!)P?����<�O�kn���3>xL�)W�ɖy%-B�0�	��wF�H���2�3�.'�=���q@ގ�d��l���[${����h3G =Y�a����0�\�`�d��e����wMy[���(��k>�(r�|�J9&�����k%���S���/�]t/N�
�����ax$��X�[b/�E@x��q��y~�x���)k~l��K�H�j�IXϫ!k�Ay��_�b#R�B����嬡3'�`Δ$rO��� n	2�Սf��T7|Rp_�^�ț9�j����e	�)1�d�|���m� f�������7gI�K6��%��jC[&�|��[!/q�� �JC��+�M��mu����+��&���أG	��Yz����fɏQb����.|�M̬��}��6�R�͖�uڸ5��8�Xed��l�UKRҲ#�$�@� �<��h�fS;<�����	
^�j��L�Z.Br����#�U��;����5�XT�ޛP�)r�	��y�;qC0��e��̪6_G���[G�ǀ���Ӽ��VJv���U�s�j�^N�h~��u �V��{�>E�؞�{@]�g
�2�^���bN5��q)A��� �v(n�(�U���wO�I�sɸ',h�<_Yy9�e�^�`��h��r�.5k�g'!��i���#�xƈau����w���]#^�mI�9�Ȓ�}lZQ>�B�tu����H��H�_݇��ә�L��x����s��!$���X�|݆�Q��^�q�&��9QD���]0/��ff�<N��D�Y%� �'�W(2�#��^�b�>�����fh���ȗr�Z��ޓ�nu=k�߫����s����siP��|�/�˥��9���G�RȚ0���ѾL �s��=���eS����ۿ���>��|�D]�d+cy232�2�6�BV�^�Ql�[L���X�>N�C\*IV�<�@�_Gn�$�\�Ǥ������� �o�٧�����1������I�x�
�t�k��`ro�L[ʩR��C�)3��Su3zp6n�@G��$H)��U6x該Y:,gR���W���`�����@��G����).�����A$Qq1φ�J���B�A�keV��� �a��+���h4��Ie��9j��j��[r�}u����\+�D�x���>qFnO�J	@�s=�� ��x|[RNI-gu����wcw<~�iJ��Y4�?�4�`��dV<N���Ɗ�pw��&��Q-�y��i�x���q���������G%ݛd�fO��Z��zi9�z`�Wo���� �(�� �W�4�V��;���T���[D�����AAa��{��{���f�]K��g��~���w�K�L�5����k��g9* ..�Q-�즞'o ��2��>0�F5'��9��Y�.���������]��7_����?Xv�ށ��`hY�_��{�?�J�,���rL���y&t��s
�3��j��I�\iu��B�����2��Z9bBuk��G}3�L�a	=�Lـ���G�p���jo\��$|�>H�� o爩��� �����sH=T%��X��כ�w��z�01�>���{��<�j��!k�Lc?L1�.L�ʝ�J�)�<���zG�#�b��,{T �ssG���#�`^�sz��ҭ���{��-%�B���z�^3s��w/UzWpp�Ԇ����]�BpH���A�3q7���}S,E����q/zR���Qb�;Y����%oI���C����փǎI\"��j�{Tn�q�@	�ͳ��\K�m�T5�D'���Y���C�0���h��cU���^TF��i�[M��x&���a�����Ý�>�׬X�:nH�N�瞎����M��Q.����KV�{PdŃ/Ӹ	�5T��nߛ
��d#w�����������u�P�:@��b�6C^�-����;��?SJ9��_��M$�	1�5O«Ȝ!�I��ř�"w��6 �����6�>���*� X�,�hs%�� U�$��$���E] P:Ճ��T�FZ��+����4�,���>*�a�s���!4e�}'��ԿJ��Q`�A*�y>�6���%��7�"_@-�:�cJ
��f���1)�Y
#��������>��<�+3{y�o;�2>&����i���ս=
P`�-�3�qh�P� �i�R�V���Ǎ�:��wD��v�9��2���#wd���ڒ=���h&�b��Ёg�=�L�k'O��Z�)�� K�Y�dWxI�M!$_��x���c̔��_��Kc2�a���lˡ�?�ڒbԂ�u3\�X�M�j&[����+��S��ގl{�����u��骧��!N�-㷙���sN�{e��� �ڢ��7�dV��/Y����!'G �=��m?��V�<�J��Ӵ
<m���ω=�������!Eg�:v->}O�u��	2`�����ďI�5��u\�U���"���H��2�7[�A9�:�U���+�|�u�6�cVmb��o'j؞;�K��5����:S��ȃ�/�����^լ-�~z[Y�k�I��gV��} �{��8O� ��`?;�cI�9G1�����/&?�`�l4���W��f�-)��ZMf��^e�!�y�58DC�'q^S'��T\v3�0���B�Z�k;���x�y5�韼�DY}�V��2�j|�+�?�Z�:փ�?& �	@s��s����Ȍ Ypg ���,�f-$1aXaWs��1>�݄�$�-�����Lk9��r] |�#�f��sM�:gUo;\�
��3�0��������5�kҿœ8�� ��A���Mc��e'KdOFB�/���s�U��Ђ�v��j�	��ǾS;��?&��xཀྵ���#�x��[W���\�r��#���~a����贑gl�
��~#���
���r]�[Pt2b��57�F�W�fs��t��X������FR=~�n9rc��N�0��Z��]]/��S믤�u���㷭�jmltl{$��śH�m�����8�9g̃.P�N��>�ܓ3O� P��F��x� Ӣ뛐\Zrq�K����]^�lDP�ڹܨ���Y�Q��I��3lh6/��׼��	*��SV�%���S���t��1ۥoa����Izp#��^���M�RHV�l§S��hHxc�ໟW^v;�0��D?y�Q��m6�2�kf�Q��{$�/�!��0��(��Z�k?�m��;�p�V�=�x����% E�g�DP�S�fo$�)���b�}܀�ۨ��u����Y���x�Zj�4uAj�������d���Y��#'�6h�,�cݜ���$DU�/݁�>F�����R�q�����][��KW��s�5����$�VI���Уm[i���
XCa�/��U�mRL�&%�^�N��'�(;��>߅�#�d���j��v��_랻ל��P\zBjx%��=��a̹�;n
2�x��/t�A�Ң��z��̿}� �� �'r[ȸ"-��j��%+�TW�6B�׌�an�W�ٗ���'�x����e��M�/�p�N2u�&���) �3q�Z�!-/v��b9q)nxXW���Վ�s��X� ���������dT�Y��?��� ��¢��5�!�R����M�J�X>�
 �x=�Z;c�f�䍙�j��-��
�E3��Bm����S�!����ͧj��߰��.�zj�'�V���z{�#^&�b��d�>qȋ��㊩��L�ΛS>]�}�F�	� X�u��i�x*���VL��������-�`���4Ot�*.S�޹�,�@�eL���V��Q���v`����E���o��7)���!.�n`�� �5�Vw/Tb��m%�����S��u6{�
��k��2�~_鄏U�x�C��=��C������D3.Y����|q�p����E$y7?�C�d�F��W�����b�?��E9�BG�l�wJ|:M�����yT��[6̫C=�o޶,�����D��s���w.L��l Owٓ�Q�`��V�7E�}��_�DO�|��j��$JJ�Bh"��_?B�����؍��[+)���KR�60e�ڙ1r��)a������⧳���R�b�˸r�3�������Qm��CO
 �rk���F{�1�V�M]_go:����������������� 2l��Hy�e�\�9���|��H�X|!c�<kV��VN<��B�p�5��MpQC�e-ҽI]� C��.70 ���_���i?+6�����-���<��j�־�\G�;���Z'xgF�Ԣ��IK�����[}���F��ڐ".����r�A졉���h�}bYX�w���p�p]f��w$[}����1	��vWߣ��;ր*��k��+�����d(�w���V��ئ�X��Uq��i��8)b�}k�BY�L"��@38��0�3t(9��1<.e�u��ʛ�0��T^V�J��,I���v�����S��H����H
k��޵D�k�#Eǐ�Do8!<p�ũ���ٵT��/I,s#_&s���<����I�.l1��� �j/Cq�ֈ���-�/t�I��?�Xm/-^릭r�Koٮ���-C��W)�)�6�H�_l���hnq�=||���Ǘ�2S����,�e�J��-p���O����\��8US��Sv�_;���O,(^Z=i�=�}��b�����".d�jt�٪�[� ��	���������y����z�J��\���'Sa������;��\7��Ȱ_%!�t�w�B���O4SM�N�� �\��9��W�HV���OM���K�\��a��ė���x��pʆ![�%�:����?d����1< T��T4��3�)ۡn�P���>5�|^�p��@⬨�4������4�3�2�~��_�˯ztn��b�n�X�F��g�����K�<�8e�F򵓚<��b��鸿��*��9��5���+���M�L���l���ݖG��G,�h�������7��#��Pw;Q9��
:Z(k��ͻ()z��c�y���䝩�T� 7y,�_x�|J��קѺ�H�ݸ����6)	����hi�2b	�,,��Fԭ�NWx�^IwV�&����*��I�֐��V��DE�����ǒ�O�^�ޭ��i���Vɗ���L_��j��oy��׌�8�����k�K���JJЙuc�j� 9Q�O�V��0B��x,����lt(��j4�$���B@]�JԞ�v���y^�EW#S[�.uW�j�%\����p��\l՚/2.|��V�wf=֚� �eG��Aǖ����6�1x��ML��u%*Ѷ�)geVe�eQ�XF�%r0��K���zi��a7~��Ϫ����6̞���w� i�Frw�L~���(e�q�7|n_��[���ɡ���e���a�Hš��,]�Æpe��kjVT ��ӈ�Ǵ�Jd���x��|֊��uUuF�v�3���c���^N�Io��S3����=�G�����C� �����t������-�X�a�"�����B�������[<g˔F�Z�%�"��/	W�e��<�g=���O���)�˗bG��DL7V�i���G8���3�h&�����}*ɞӧs�]�ItA���,�����he�3~�r�>7����Z7��.o��Pm��j��UҪ�*Zp����O�Ӿ���y�v��cI64H�g�e`����F�LC�Փ
Êн"_]�W���I�j��4��j5(���}��S{��̙Tsl�����r�$�C=���+4�,RF%~�g����:,�uR�MHjҖL$�ڐOV��G�Z�76J���-�l�[e�c�l��f�j�����5ˉ\�[4<���y�t]��Ë5!�$r��ߥqw�
$��щ��]� �!y&�����Xl����V�B�ن�����;�B��\����yA����i��v�T��xGz�:�$@�(3�,���GV>w�FXk��� �瑮Y�-ѻ�B����ڶ�J���]F��k[��K��a%�t܍�B��D��,4"�r5��K�G�:k�P�cU������X:.�;O�ט
ڒ���a�����~<fbA��X[�w4��`���&Q�O���l����H.g��^5��?p�w=)��vU������}��*]t���_O�I����d7���VK�q��	G&�}�����eJ�3N�x[�Ζ�A�<fe��R�2���r�5�s�����d�-��DI�T6P袣JYբ��fIz�����r�rz(?�wE�������C�W v����l�W� �n��M&
����҅���Y%��>9�)��㮪�wx;g����ȷ��}�����a��M���ಊq/�����8���o�ļ�g��q5������^W�i�T�̆ њ*Y�Mp�?�x�aXb�3�ho:ju�=�C�ʲ}߬k�e�"7g��t�C�3�4��'Μ�)���Mo�鴡��7�@٭��u������l�f�C���mr��ӥeÚ���w&+��k;�7�yM6fn�O�_�4�i�/��_�1G����/�@w�xa�7���)�u��f��|G��y�%U�np�L�k+���~/ؿ���=3�8.;����+qI��a	ʻ��KQ��$��Z�1YM��}��×N2�u5O�L�_�ļ�J�w����-_�ua��$�\l(+�LT������+�cmQ�"�M0��ђ�1)��h;7�o���$�?�@�E@�4)����?	Ku�ϖ��Q��;�Z\ibW���sV{�)�C��`�X��M\	���zM���r^`��;Pkȴ'�r#W���).������5�'�T��\�7_��Wh�J7OGdK�Y�ȮᕨY��X9����	I�Z�aiSF�Rړ���]��s�F�&��B#t������k+xj�A\(l��>�JEe>K�w�DQ�����M�yo�������/Lk�֌���?����ؑM�Ԙ:]sӏۖ��Y�ܽN�E�����C���]�����G����\�
7�MǇ��,�8�ȟa���a�ݬrt�j�rJ�/�8)M5����C�=V�0�(��X���ߞ�.U"/V��tV�C��=��H׊�0�N"Bdsja0�+ETX���.�Q5i��°�v�ˋ��ߒSe_�\�g]Y妛M93��9��់`�B1Ӎ/])��|�+LT)�m����E(F�X�<f�B�c��KB����(���n>,!Ry��P�
�
dH���f�i�~R����d9X��A!'��*vR&д(&�Q��U�to*D�<+�<�W���)%�h%,����ܻ��}F#;���Ĥ� 	Uc���Y��Q�����@��Zv����usb���cw�b5�PW�Tz]X@#� ���r����T=��Z�,��j�9MF�}�+�xe��ӵc��/J��\�QW/�2_�l�c����U�+jXh �i�ݵ�����%l�vW5VN�zg��	���1��N6�? �
����P��dǲ���c�62���Q�F�X]B�|�F�G\-W�5�`�V��a5X�p�p'J�~�*�bإX�֔M	���{*D�-�Lߗ���5���i6��e������g��q��0%ɡ#\�����ٓj���F�Zl���U��f (y3�2'��Պ����_6\}�#�Nѡ�ϙy�F	Q4.t�Ӧ��Fp����c_bɗ��3K��k�ZЂ��o@�
s��^ۖb����e�K��H�0(��;�8������T�u�#/��޾HS��[�f���0��'բ\̓Sǿ:��ػ�M[��X/�O�Y}d�ٓ~��̕y?���C�bV�@>x�ι ���%��c�z�~A�>>O���Қ1�.忒�o����P}��Jl�{}ե�jp-����D Sx�C����>�t�U��`���z�Z�_�+��� �󪳩Be4��\��ol�|Oʞ�ܧz���/#f����K58��!Z��^ᤑ������~��h���K�@��υ���!�������˧��E$&}��FM��y�\�x3jnݲf~ej�V汀t-��>�}����P��M�77�S_7}�3* �ؕ�����7�q���v�/��H��%~7���ԅ�90�.n�:c�ds	VAM�L>Ɓ��Ŵ3����sunof}x=��J���1I)����+l0���"�O�P��/.�$�^5����<� ��ȳ���`��Ԧ./6��eL���i����ơ��.͔8�f!���x�Y�a�n�>�SFy�����N�������L�|��&��'���c_�6 �&�k1�pև���a�KⒶ��+�kr 8�*9t$�BP��^"@�)<�{>�������Q@Gɗ/�D����a�$ �y�Bs�A����ᯟ�-K�}&_E���������Hχ	_�n�q�'�B���B������濾]�\S���7v��(6,o�H-X�{�	t���͵�ؔ�t���d&���c�A� Jiͨ�ɗ*^�>��[yI1���4�D E'�����ڔ2Ta+�R�L���Kf����̣�4�1����nh?���a	\wF,v���8Bd�ˁq�y~׋�/ {�7�M!M�	,lJ�Ǽq����s��H�g����C�yx}1tMS@�.��!U��/W�ڃ"SR+hqh^;���/����ӕP�5GgE=���Ի`ݒ��v��t��"�c"�51OB�&`��/������йu����L�rxWΑ��/CgӄC����MX��i�%�?Xw��xj�w�j�t�-n��.	̒+/�Q.�'瑌E����o�
�Yq#�B��xy~�0�� yn�g΀�PQ���X�{��L7XT]R�e� ]:�E� ���ڞ�&�+���H3kVX����/�
��iBO �oS>&��><�rL%g�-�{�݄m
�n�7ۼ�4VK|&v�W������3��;0}����V�F��^����ӛ��i���7}0F0d�=_E&@��7ł�,]�]��lH��\Ј��(b��b��f�+��;w�Z��J�D��i�m$=��s̑Q�C���yh�}N��'�����c���C� | �	eA�����ε���tǖ���"�ڴ{]��V}��O#>Ȉ A*��x�U\Q�q���+������J�a�-����nғXuZf���스1Cmxh9�����jL@*�)�����&�(o^���5��4�U�:��DKu�g��`3{�Hf���q ~��B����|��P��*�rW��R�S>��O�k?���D�1~�v�������<!;�f�9x�^�nG��c��)�C�Q��e�P���|����T ?��m�h��$�|��s�ϒVkމ4�,�]�Eс_2=߷B�~뫄N熫~�c��*Jv;6E�;�Q��9ru�c�.i��DG�>�oJ�_	V�FҚ�3y �:�p�>�-��G�80X��)�>�\}}��r����jw�|����K ��7:'B�4�N��0��b���C��2�Es_$��Ze�
cO�f�:�;���Nl;9?K�1���Fs�l��>V-�!����L�a��,@,�vN���ɝ-�N���mcGF�\��r*X���n�[�<F�'�%-P�9��[[��[�@5Y��d�Ł]f���>ǵ���оB�����؇�%F^�t�&�)1]ܐM�*4Rw���X��t���S���S�#����?�o
����{����^��k���`�m-'�d��_
md�`RJ1�.<�<^���R@�Vm�vБ�1�!�F�#���M���uYN �E�����	����tj_1�:f�KS��iW�Α����_�BXN���A^1)+�ޅ-�?d��<����i�2T���)اί�����6��yR��7��3Z
�9�	�5x9i�J�8.@�d�L���|rʐ%�G����O��iZ���^a�0i�:|ްt��/*�;c��[�"tT ���/J�����Y�@H���+=�<ŨMm�@75aͅ��
�i
��M.`�SjSٚ�q��8�n����Zz����y�Ou�t�H��'�&�B��a���d%��A�5 E򿩿	1�N�Q]��ҕ�dͲ��<���{FV����22<("�\�hH��_�ȋ�L���.���,撿=d;�.U�&N�I�	��R���eTw������D��M�,���w��ĵp��[���/� ��-@Ҝ,���(d�r��>���mc;Kv�Q��3=�J�)@B�h6>��C�/l�a�OC�jpv_�J�A���?S��C�YC�:JP@���T;���2�~����s�0�S�+J�����֥�.wVU)�q�=���7w�1�Ώ7[��1a�Γ׎=a�<���g��!�V3k�c[��c�7�Y�;Ĩʦ�偩%̏�,����$���ԇ^FQ�$)yV���e�����g.��\h�V�߾���d�KS�.�i��w �X�lb!U�R�1l#��ݺQ�ݬ���=%����s�F��ܣ����s�F�P˔�k��=֬��ϭ6�G��4
�h��5��B���� ߔ.w�!�[X���MN�S���iG:�I�p��`�cn�݂$g0
���������5�$���E�$�&���D%��К拿s�& w���5*��j�-�K��J����G�RҒx���O���H�!$X�I��t��h/����}���k�fژ����)����Cc�i²���� �߯f�!ȵ���ݱ����]����Gj%�5:�ix�������gC����6.�dZ��~�x�2E.�T,��Uep���/7oH�!�tf��T9z�N�=/.L-���F��|x�he�i�ӎ�T��\rK��L�狳�5�M_ą�^$ؓ�.Gy���=/�W.,������w�������b�K�:�Ug&k�ok�Xfn�Y(��Ӳa����
��+c�X��:�6:w���p�E�b̢��w��Lŷq-fZ�vn�>J@��2@}�	�4m�Η�@�����;oD)�1Ԏ�O�P��?�ک�5Zd`�Y�-�K��������*a)RA١������:�o��=�O�3n��5�&�vh�ٕ<��-o��G#L��8 %sљT�Ցu*���z��O��+��(�r��Vq%�i��#p��f�_4�wn��� ��p�c�c&��:� AP( K9p�����a]�	�1a9#�ze&s�
!S��}��eP�����4T\\�jťƤ�>�Ǳ�b�,/-Hp@Z*�$�;�m$�����՗����j5�};�������u�F���[��4�lz�O��e�c����	�D � �^�l���jG?���!��+ݼ�z�R4���|$E*��@��W$U5*|󿭺�Ӣ�V��;/�NN��y")P�����dCԄ�*bF�����j��,-���8_�������^Yf�O����!��1�rX.�xo��'(Z��Bi��Z;�G"'޵R㺋&|��m,�I|QO�f2i(}쏕b<�oy_� ��@���i/��IPL�̥r��x%�)��k��U��R�]Ԝ��i4���b�e�@�ha(�}P%���CH,�\����J*v�.�
����4�j��Ƽ���4۳ϳWͨ�UĨ)Y��r�[W����0p�*���*��6be���@k��Ƌ��G��t��(8s�kզN6ן	��rW���jX�j������@�r+�^�qu��$y�����������i�UNm�GN�ú�E����F�ԕ�ǦC�T�v	Y�	�}�ݢ�і=�7F��?t���l�pk�g��<F��]O���v��> �N���@�-��|,T���:Ƀ-�4��w��a���/�v���J5����y�Lg���_?�,_d�d�VP�ü����ĮM-��LW!E����)B��#�Up�M�i9t����lI,-��k��T��t\92�g	0�i��*�dÃ�-ZU������FW{�;�%sX9j�腺����YR�>	o��m�9ɬ���E`�4e���(�x��%地`���G�!	\T9yv����!?�M]�������\{f�*Yj1�Ez���r���h[��&�$^��fG۱�y�Q���ǫ���xh��U1����X�Α�wm���7	�w,���ܧN�|E��Gy�s�2j�V6���/��kk��t�;C�6S�]���3G뺼i՝�T�j�.)����0�5�|B����Q)��y��V۫��H��ȾUZh+{]Z�Hǣ�T�R�\F<��t�I��M�흥��Y�;��XY�5��ۮ������yq��c���ZkX�K��<�5�]�n��� �$�`�G���Q	'�ms�=���H�S��*��p�!���c �Q��h��j���f���y�U�ֱ�;C��ڍm���V��jW�+����'ᵛL9�ڧQ���ŀpY?��[��
�o>>��un��7�c��>�]2/���LǗ��re��R�iRD��uk&���%��qY�s�&Y�����������%�<�����$�T��XM���l ��ګ	vړ⺸o���{T5�\.�6g�-�A�_��|��B� ش�h�'�Y��O�� SZƨ�@�M��f-.��[W����O���a�����2_F)�~}�����ܹĺ�b Yv������k�0���r��c;�vm�$��)������hn:E���xT�y� e,��?�[W�H��:M'����a�B������SH�{�.s�fEީ�IA�<�`z����ax��d\��%m[�KA_��m �pQ�>ƺ䓈H�D�:���R�|k�j)���YKk�ݨ�Z�Z F�+QpfGX��7�X�6v�9o�hP汍W�Vx&^�%}�f��-�<��>p���B.��?}pQ (B��kP��m^����B��x��!0�ѫ6�x��_�h�w��L��f����a<Jfl�~���w��ٲ@�1��z�!A��A��O�y��!��v(�"<�� �����c�̗�b�(��	:�c����}4��:u�Vĭ{O�%.PW�o����Xb
$:8t9,r5�;�L���P?��H��c��Ee��{c���T����"ڜq�,����敐���s�0�Bn����)��'����2�gk��>oV����B6��"?K�8�7�AY���Cא���S�nG�඘���V���^ѷXϴ��\Oq��RSb6��X���������)\�
}�Έ��r�����X1��/�����G��4w5�v8���k̜�`婛�Ƥ�����2��⼹$t1;�B8)T᪷�]��6gE|F�� ͂���G�k �$D�TE���X�N���#�ׅ������F�C���_��,_��2zi�#�Sh�?)����a�&b���Z��sU�ێ�a�d6G��0�|��J8	hG��Pu.<Џ~Q���"�u��TpW�L�x��Ȃ
�i�`�-8/�}s>_�^��U�i	��6*uNYi�-����\����w+�Yw PT\�������|���]��l�߅�hi�&�Ŧ;�ݟ3�\\�3�{W��C���m�ѩ�wD���"_P�)l��T?/uT	�"Bvj��"V��pv���ts�vk�#��C�����b��ܹ��z�����܄m��яg1�?#Lrd����Q>�Ypw�r6'�5D��w��Җ����
�,�;i���O�3qԤZ�ᓦZ#�C�q������:����/�n������Ғ-��7"��� ��t�D�q3�o���	���[uoP�]��E~�����z5ռ٭g嶓(��k�^&%��VG;i��p�8�ؿ�k#M���N%���㦲�'� J2�Xa��Hn��[V���J��搣*�����!�\��`\���:Y����5�
�����t#�%��J@e��r��d��}���]7���YiU�	d+��0i1V���\����s*��5�O�?��p�B�\۴q�jWV�����j��3���?�սC�o�_����'�[��؉$�ܖb!#�����顰^�<-L�s�Nʎm��m��ݵ�T��ǲ�''�;g�4x�ۡ�L�l�"�:@�J����6�N��@��P�������<O�Bk��gm�tm�a�Kn�f�m���r���>}GVC�}�JD�f�d�P��$g��\����+o#��<x\?0���|6�vј���ުަmb�$�)Γ���Z�vJ����]�Y� ^v�,�2R����q�"k�E���I��P���>����0����9[�lH|z-�
̬��@^�	��r=���K�Ŝ%3��\���*����@���+6=br�3�W�k��%�������L��`ak2ׄ��!�	�-���lHQ<?�Ɋ�o6��� p@Gu���_��B������#�W�U�:�YG�خ}���|2km6u~ۛ��ܟrR6�N6��SL�!�r��t�8�AN�����=�g�8��h� �ɾc����9
)�C��§��l���'��ە����PÃqV�o�E����ݧ}	$�&�>���o�<��]�dP�V�!Q�!`���*�Y�l�uɀ�I�uq�nn����5���w�K��I˨C�]?��`�%�G�6����!D�E��t^�z_�=Vɘ�m�3��g&�3�f���������������C��Sg���t���0��1}QG��0c��XX���d��� ��Ѣm_��ˑ����'�u�i���&`~��=D�?���涋�� y��ohgQ,ԡ��g��������}
m<~��.R�n�Ԓܒ�n�2�6�_��6�m�����h��X���QG��}&v{�^7���浓�T�L��K.�VL�ݹ����
E�!��k}�s��o�b�Xb��	~�ɨqk�b1ц��7�ɓ"^e��H��ƶ1�-�Ҥ�SE�a����< �%�LW�Qk1�D±XRP�{Y2�����~E����D(I`oi�����)]"���Z^c����_nF�����r������/������T��v�#�aʁ��ҷ��UwsG'��eT���<g�at�.��5���HxN���,L�d�
*�� �.v5�>����K֛I����m�R��
 �72��l�D��	6vSGe�f9����W�*S1�X��Z���q�oV.V˖�?�&�q��b��+:^��Q9�(D�[���Ϳ�r�;,e��%vh����RM�^�i����l�:��*�0"q�RX�	�zp�N?d0�e&mxG�a�۬��>�o�#�F��a�q�CZ6��t�h�m<�︋�d%_���&P���}���k�.�s�_A��?���ݱI�"N���'�?�	�tx1)+;)k33='�UG=�܆�c	����pnx !4�F���bg�Y�/�V�6�U��u�?7��lcG�*O(!k.5&�q�����9�\ZLI��N&�.�	�89�L6V>�˖���䨩(X�H�C���O���rɣkWd�X��i+M�K��N�f����ʩ�hw~Vo�kh<�(�����'s�GMea�nP�.^[[�$i�o�Ts�������.��m���_�Q�&��z|h@�%�c�v����0�5>��s=�!�⹡X*�$Ӡ���Q���e�v:������۱���BO��|>�~/���1�������(5{��g�l�_l���?�WB�n���9�5Pe�C�ǒ�}%���=��"C�(UzU[!�C��g\�t���f�d>oж+��Œ��&sl��:
{�]�,�W��f{�V=I`��3�` �l���-���j���h�2l�n76�ߧ��:p���d�υ�s6�q�Y��p��<�g䚕鵼7{|���MX@f��6��qr�����`�|?���>����Ә�?�O���)�E�"[��Dɧ�<�$�\��>� ��"�J9���.�o��)oZ���;PyЄ�F�7Zn~s���>��;��8Yf���;��uO��}o� 
&�q�ޑi�kO"�� |�SR�M��i;k/u9�.Z�
�+S���� ����r���~}��2Ci0���
����e��f��Nq$�pf�$�J�!ҳ\N�6���Ra�5���|S�U$�~�� 1�C)�����2|��]�%���R9SU���?ơ����lxr\�7�d��]/��_�����38�6*?6��P���8�xE�f�8w	��Rt_��\O�o�`H��x%D�b�p��7H�}V���R�p�C�r?-��[��.p�M?�)�Kr���d.[#5RnLԃ-v��8l��?\v�}Ab��B��k�כF����wG�"���4�TU(d�]&÷Q��WV> �,AT�;?{����\#3T������*nGa�4�L��UĚ8��E��bu��dՕ�4q}��*�W����[��
w�3$9I Pw*l3&$Db�д��YQ������PUM'M�	>�d�T��N������ڍ家�m�vZU|��h��k��������s6�@�0�v�k�(�� y�c����/X��mS�T`��O����~�כX�K��H<��H��i�*��i�(�i����M��'UnJv���#w e�{�Y�5�|j�����n�2��efL��ܟ_�]��o��N�q��H��u��IuH�_��|�݁�*�1n��iI��q!hu��ct��W�l[�s`��������[�гJ�=\�4�T�-AA�G�I`�[�����~�2`�"��N	�F5+b#`]>`�+��(^4;�Y�d���b��ee�v/'�3n�gms5���B����l����qN��lﯲ\��wUsu��@�K���	}9�Q���(�X���1�s�3�޾:����,㟿}Q�XE�w�^i�������6[���<�6�|sl��UCn�+t�����y�(w͙ctP����������?�F�Fw�"��Ϩ�?� %�
FWs���z��Y��[��:��/ʵf<8�ϱaկ!C�h>�4��T����*��N�1�U�J�c%�8T*w&b?~�����?�@݂O|�r�V��h�qNO�x���v�����朰}\�J)��Pܥ�e��Y�I��|�����B�i�x"d�z�w�gb�QN���q�5�4D����	�M�um>��~gTQ$ӆ�L�K }�,�=�5̏�UM�~�;�7ͳH�[2���U�S�3�}gݒre?�O+����aH2��-E���@¿y?_e!����~$,��5);�7w'�4X�\��:�t�S��(}���"e;I�,�t����咵�/��XzU.y�n:8�V�6�۳��V)0�6���K\�μ�H<��P��#A�PT��v�0�����s��c�^�@����_j��{��{��P��}�<���x�ap�>�ff�ӏA��4��Eë9=��;��Z�@��a�@���U����/xBy�T�f�������	? ���H.�_�u�[Z�ǜ�'\�V��:o)�WEW��uD�wi����΍&͂�v�ro�bP�G�)`�Ԯj|kc��svDu�u�<E��K5'lE�OՓ�T�����F�g��@�(�p��/�C����ԏ���]�Ӳ�	e����g�i�2p�|�"Vᓂ^��t���b�]��D�)1w�h�U?;�?�Y��VJ$`�v��}�U�����7WUe�dm�R�%�秂T��w�ԙ!�z�1or�����-��0�lC� 9�UW�|6��ǚ��@��DF��Y4��6���WQ����>0k^�5hK.J�>jw�]B�Nю�>�f?���z����<zG�5�F��M���4�߈}�_���ztz5~���+��CF��� e\z0�}�\�m\��e,��$9̏�s��_ۍ�h���=y-7�h߶��9w.��d�f��v,g�����;>����;��w~@�|���eo��+�sgq�9���*��&K${���e�4��C��������[�~�s�l�h�1����i6�#�o�:����.�{!�����`�[�!��xc�	�>��׳�	T+2}�1i<j>[z>�(I,������<
����Z�����79˟-��pw���/�p5_���ӆ�-���P�}�_k��Q��j5xЍ_"��T�1�T�b����*ϑhX�"����W-��{�ݿ�%Z� �41��;A�� �Pa[1Mw�DN��Ơ��i:�ru�%�}��<�a��<홇	���.̔���s%���������P� �My�����3�0�,��&s>��s�D�y�[��o V�����0���]����O��H��
��~gwf���4�dB�7�zq���@6�CY��]�#	{J���Yު��gO�k���;��O��{P�_	yj�E�ݩ8iT����{4���y����whg�XAR�s��s�@�˧�ssC��:���k��āF|�������
�(CT��HC_J����缇�^��k� ��;�7�o[,n�詘�ǈt?�aq�n"V�74C��*m`���a�������̰���0�m��9�q��?��;��r��'��y8j�X$^��@��b�9*��k.�f�3,��۵+>>SH���_l Rt�9w\�%rl�p�ju���Q�Y����g��j×�i����Y����p�ƴ[�Y1w����v1um.�pI���Eԫ�2�o��q�E3ī��D   5>���rl ��brY����Kt����ϥ���(U_R�rc��w�;<	e`�#�����3�E>����5�*�M6i�n���t�d����O�Nq�غ�@��3�&.��U�6��3�����x�.���� 9�E�^|Y�9^�>׺:�_�#��&b:˥����S�QByu�C�R�*B�����ziۄt.)� ���K���  ��t��tI# 
,JI)!�" ]"ݱ4�����y���qTv������ra
R���z}�/Tӑe��N�#�[o�ֿ||����١���?��z�zWd1b�Ջ�@�wK�t=�Ë���%ڃ�i�f	d����UN;���׼���.¬.V|>
v�;���~�>~�6-^��۪�0�,��޷���T��E4��}־<���6l�,��M�d�\�����W΂��29ml�[�g7fO�v��
*�N麭e2O}���_\��:��Ѻ�a��
=��7 ����`�|i�Q̶�+��`����ۻbf����{�~����"�{� ���K�$�.B����jXw4�:YY��)�tͲ��z3�Uj,��m��qz�%"�֗��x�V9&��"�To2� ;���d�YB"��PV���ɠU�h�=�F�lim���0])\�u�� �gZz�J�X����������n��^
���g�?kZץvͬ������
՛��<~F��^_�g�͟��[~�n��lQ�%u�������,��N��VE����w��˽������??�5�z�X�BK���w`�ef�g[���G���S�O�T��n]�F��h���ZMa����8���b�*=���r )��Qs��ec}ƾ�O�0���J�����2��)�`7�obg�W�Λܞ�~�I�O ����gn��r�x�ԡgg��CZ��*�o1˸|�+�V�XN8s�歘��7�S�E7H>Ov8Ϡ8�qHJ���5���Cv�8J=.��b˔1�fE�H��v�k/w��>,���Ŧ�8Q���0�F��Z�:��t=n�^7^��o.,F1�g ��y~�m���Bj.'g�|��>�+wR%8R��Ij0I�1�_np ��2��{4@����+
�	ؿ5�F�����[?�Ia�"��{TS4��fi���ٌ�ź@�j�ﲖ�݃󲻔t�U��NuIW�����C��$�/6F=c<��H0L��9+�1Ҫ�M��e�*��Z��.�d��O�RV�|�'|~�)�S����X�+���	�A�@�7t�h�g�G�團�����d� �t��^�nx3_�׽ay���е6����̴�����n�@���������,܅��,�r��%��� �a�6e7������s�#����Q�������=��7�hhU-�/z0���1����t*�y��7"�?rdU�
6%lʰ�I��㺎���]�e<p�¬T塾�����<ݮ
l�3?����yt��B���{�zoͮ�s��b�HDW�A�t��"�G˼���^^�hZR���5���/!����R���&��tF�v� ��d�%��?��u�T��R�s�g���WA#����~1P� K�h�����SB�xt���s)p#��"\���[�ܺ_u8F+ȁ����W���������vy����Xp4���lQR�����g�}/2�^9k�b�7�5���y� ��TR���~�oט���E�V��%���О���S߯�����o��o(.��P�:��L~�ӣ}���{Ճ`~v�_�S�O��\׮��Y�屼�qxa�q!���Q��ηッ�S�'�����ϐ7����{��)ݼ����)��*/��}A 5�###yi"���O�444�w�il10�K�J�G�G.�tl�I޿%$iH�A��$a�w�I�gB�M�e�9Z+T�X�ⅱ
Sf�x���~�=j��.s�U�����t�������㷪㈴��{�t�!��R�t�So/�O�Tp$w']N�|�G�1����W#���$C����ŀ����ME�WS����G�|�Y�[�<��}������FG�vww[��+���:G�z�A�°�T���=�����,��`�q)�u���U�t&����ۇ�(ޒ? ����&����4��#2*Wm��j
�WW�pt���)ьx�w^��W�&��o>��*��W��7�1�#�AlY��_0����&'��+J�[[O;:X�M���e�,֘[��n��se�Q	b(�
G����Ì�V��U��ߊk�g�A=�[Ε�1���ѺS4���p�0���K<N�������;��ۿ�ONm���\�jE���O�X2޸�B��@y�hz[|������f-G�^\\�����>���䖐��*Mnmi�655�'"�9��)����h��U���$$"�����{�X���M܄��N�J���l6�}	������y㱆�m��7^޵�M.z=W�^���^]�ϋ�[�%F�B��&��ţ���YG�2Ҋ�R>���;���J/��e�~\6���.�?'�-ύ��8��f��~b*��)vt��9�+Y��6�@��B�9��c���KH0455���I3G�LK�LJ�00�j��R���aT44�-�0M�����\�������Jh+*_��_�3V� ��e�S޺X{ځ��] �[#ܜ
��� ��q��*d!$(<��{v����G����v>4$&�㠎�݈�ř6b�K��y�R�e��Ku"G�'�4/[�m�e[���x7+�)���������?⇇݉5*RD"O��B
�	��d��o<��CYW�?�������F�Y�BfV�tth���g77�H�^�����o��E�B
;�m�����ĞO4�4�n�گ��nѧs���X��>VbR~Zy�'�w�A��%�46]1��W��JKgk��i�XX����|��qyz�:��Bj;���{��b��&��R�#-�aq���w}�=K۫?�W���-��q�C�-C8cdFG���(�^��������Y����*VNN���öJ������Ӏ����tq{�fw�;a\b�`���1#Af��8K�����ȯwX�[���8I��c*XM���R�g�1��ѝ�P�c��
fI#Vm����Y��-�F>B�k/E��ju`�c2�7���7�Kte������Ӈ��6�8�ﱮ3I5��H=�&���@tgq�3J	�������F}V��h|^�")ɨk���z���g�acoo�g�ںI���g�d�$Ȩ��Y��VV�)��k�C�&�AR�6�������:Z�->��SG/&�dD'�
�������X}�`e$A5"�oh�y�~�|�Bi��e�K��9+��uLp�e^��ܗ�/�H&�xܵy1��MS�Kn5������/Ok:Q�2�Cvv~�]
*��|(t�����H�_�k̎e����C."m�0Jw�33@M"v'��X�s�#�nh׾�#+\X���l�l��}��r�3}�N�:���sN����܍/���sh�fvUE�k@{(�
�y{e#q��9(Y�7~`��e�ⓐȃ>���1royt|��KGDD�&'��a��w�?�1��u��vT@CC��3x^J�G�(�єOC�_O�M�����^O�9��P�"��(Φ,��7�>m1�&�T�2�H�-1���R�K����D�z��z�;�����ֿ�^��#q3�S�,nC��(:���Ë�`��B.���F�o���Q*y+�0���~%U��)))HX'��1�2Vlc�j�}X ������x%{��ܢttg��ӄ�W�]�.a:
�C�<.)���ǳ9���o��}�~\�;���{���U�)�or�O±��z'���Z-A�Ji֛ݨ�-)`V_>�L�qy�ĥB11��$�����E�q�`��a��QE�	������xx�u|����꺀9�����}��o�V$��a���u5����e=O`���	�^�oa�V��+�HY��,��p��%=�p��O2^�ޠԂ`Fs�ʸ �|d��2�bϟ�H��-q��e��*�?[u��ݡ��KSR1��"��� �?w�8Q��`q
N��0�d��9j���C�{��DFFF`��T����]w�u��n��rYI����wж�� �&��f
9���~-U�������Mj����D����̙MF��}2F��1���z)��ܻ'3Kn�t`<'����f�]�@�Ysu�DH�}3�b2����O��/_�̸��{^ߐ�0��:�Dx;	��ݕtOI]}�����Ų���/�{C�V����m
����}���i�-b�q�^5~ZnS��Û0�:���ӝZY�&K VԒ�����@��b�w��S.�6�~��ш>UW��x� }�@X.�H����u���t�S�H��b��z�7��ha41";:�����"	k��<:� h	�oj4��"&F���`��0}ą,9n>MZ�/�=�ߺ%���,�	� ڣ��V���O���&�1�(~s����)��m?���R���X߸{�g?���������ނv�H\�>� }A�D���iP��6�Yמ�uX"��[muz�pE86�F����
(?���`b�BLxq~�28��o���:ܼ.�)$���۰���n�ET|O��mŻ.jh��y3,�[o�V��N�J��x.��X��a�x$���y����a��ک��F8�,3 8��zkvnQ���SjbJm!�+=CB	����|�ԇ����@qc�t�+Q3hf���V��Xؓ�����!ܴ%��y��r�������Ջ��sݶ ��&U_��"����������t��q��%�k��d'N㞱7e)�Y&���_t����t���X�7�LN*>����� u� �U�~��$K(<S�c��[�@ x� (�nU��&4�&L��4q��5{[g�����G�SI�1<�Jʸ��T8<<<W;=7W9�~Ǵ=����ݿ��N�06Q�E>���&��ѝ�`�=� _p4j�I�7���瘘��Ƒ�q�M��B�&��¶ߏ�V��;h�~K9�W�,�Ķ��N��BhȿdL�tk��$�X�%������P.[���B�>u?�o{�/*u�0��R�+���+~�jOA,��	�5�0������򚱩�Q��
������0%m�߷�V��)u(7E�S�W� 	��$�rq#�f6�cꋯ-R��mG?�Wz� >9O[���6q�A�s;R_q��CѠU��2��Kė-�-�G�m���R����6�,��0m���z���*�j>��nl �,�@�:�����D���deeĆHqR�2�Eީ�gbbHcgYXBfv���\{�~��3��1�ʧ$V��H���9j���!�+|������v��G'������bᐄ��|U��u��Qc|ͅ��>�(M��=<?�C�tG��!���_QۛI��ԏ�L�k����Z7����Rl��*XAz�r*))�.�|���2�3��.ls
s�N4������6g�f�c}�P\��F���G�1�o�����/��<�|!)���3��� r����佤�G�8|�!9��'��$&j��qdqN��rX8<V+�Bʀ��q�#	���v!���H��&���϶��LO�C�U�Ԙ�4�wu7�����Y��	��S����]�/l��ߖ%�$���-�.�Z���ub�W6��9�; ����d���p��uG4�z�Y��T�8�]���hۘ�����I���xxnx�_�Z�5.�o̎��5��J?�(4b�Y�4�Og�����=�"��_�g�G��}k�bYNNNץ�E��_����r��f���±uR%J4�h�<L3*
j(
E���M<�k3�����>�{�	-Y!؝wz���f�M�����j�%^�<��j���I�oe���o�K�vxԶ��(�,K@C�ihhڳ[��n�e	��'��#��m��qP��/�@?�JA��u^P�(����<_�KWRSKP;.�!�#�潎%Nod�;J���a�%s[Cπ����Ų��<���l��P��A�oA�hR1>.��>�{a���9�Ϙ�7Ȥ�OE�0�2��蠩�#HyZ�).Ge�f���W���<Ze���c�L�~9��x����nj߰�G J���TY�?��ͷ�?�EX��c��0�q��*-���"����kC����/�:��D�B�7Q�u� �"L��ʦ�R�<����:�k��躒ٙ�'Km���?����g͇q�a-�F���?}^C����9K����ab�'o���Ĺ1 �k84�̩MnW�Y�-d����f��֔ɨ޻�����f����+}�-�d�?~D�4kV�}W�7�,��9��j���S�0N7X�t�+��;9�5L�<8���$A���u�����ҙ�SF�t�A�x�����:u%��-��&wȡE�$T3�H���-T��6�as&�=��� �[�[�>n��,ȣ'�nm���X�p}�k���Z�b���ТSv�bK� �5��S{�|`�P�e<�^d����w�0A�/
$�m`г�����#Ҹ��4ג��`"&H�|���g&��YZ����JTn�g̫�i��X��2i���(졜ު	�i�ml/A� N<b�x�p�I+c�bB6F�UB�,9`������E��M�m||�VXؘAscCc� �]`���9� #��ѧ�����6+uڊ'��|���W^������%g�]41�q�q䡲�}$�H��:i�9�yG}`��2T�=z�So��?�}��qJ�6�L	�*kJ�p�[y�&Z�q
�d�UZ��r�J��(	���hR����$�ޞG7!'葏T�W4�Lm����E�U�g&�pX�V\��X��� ��Zi��3H*bQ������8b�v��0^��;�je0Pj�Eo{�kc�N�q�4>�I�K�y�>?y𦝰��笿�V��N2����<gc3������]Bs]Y2�(�MD�~DƧg�+#E�Hx�A�;�g��uXn7�st���.�� wqJ��]����R�1Ӳ1ǌ/:p��߶Q��n����v��B�"��y�j��x<�ʥ<�{�t|*	�5�g-֡T��{�g7����yF��C������_N��ҐZ���7r��&�Q��Z�t����z���	�d>|X��5I(V��bI�$q��~B��y��\^���Bb��z�n(��)̇ZF����}�I���>	�'��hC~�lA�i���Dw�1���WUŖ:����Z�4���h�M)�w�J93�2�!O\�'u�]Ƶ�{5z;�#��2=� �w���8SipS�]$��p8���ӧ����0"[�Z��s@�X�Qܩ��gv�~t�Q����1%����a]:��V�hZ���H�W��gv,�*�"&�F(tH&�)��ҼܝH�6k�$H���1��%ht���^b'�ثX �6#���=���ܷZɺ�2U�����z�pe&i1��S�Ŭ��"Urb�v�ٙi
�Ew��9�A� .�ؤ�P��܋��1r��Dh�N$�|�H��:
���=������� �j�/��Ic{00l'<��0���D�8�q��ﮬ�v�:��I�I�ɻZ�Ab\Lˊi���i�G�p���<)�oę?�Ԛ-�Lt��J����AM,D��}�j�"84����~k,���p�|3,�Ml�"|@����}"2��� /��IH����je�=�;�' X�l�V��3�Sr��H^���=H4�m����S�8�,mx�~ t
.b��g^��	Z��s�hth�¬�p�c��B��������4�v�ʮ��<��gl8�?�a��}O�|��j��K�MAx-���@�Ϟeְ6
�E}���6�\���]Dһ��N��|�#K��u�?�H3��?��G�<B��e���R����*N�B�b)�E���I9�x[jH�,������'E9�Gl��1|"�q�zI��o���F�&�ȟ<͏�ؿ���۫�� >4f}�� ����ײA�M��/f��~�Ԣ+)��?z(��K��ZZsb��C�C��諓��]M����|.^���.�e�s�x�~�/��� I����F�"��?�*%ǉf �Qi�+s�`EΜ�w2ӂ{>���9�Ւ�&��C
��-�Q9��*_����]`_�{!s�5����ك�0|4U���T���N�5�Z��ftaf���V�K�p �@�ĉ�U#�)�ںM�`���r�{2#�Աhnf�=�K$70�������A�ժiu�Z>G��W��'�������F�%+���������J�eJ��{�0��yH��(7^ML�W�ePh�'7H�q63��pM*l\b�/����V����/f������*�� ��t�u�����Me����8�ړ�\v]�^�-�zc�͇A9�,�D�����9y<'@��V��7ExPO �}�~���4���Z����	p��Eq'������7����S�[KAg�,5���^3�gn+��_<X�Y��#z�0$a�p�a�����e^XX���@ �^��i�T�g>�"i_mA�����ģ�~fc���/���JZp�j`�������Ц��=R�.g��ۻ�!�ܸ���-��,32����E���� �=2�<D�!T(&CI��4�[�1	fsC��yv���û���[~�f	�5i��DQ�ښ�;a=|7o^;?=\&y��̻�Ăd<uGGi�l+%�ĳ IXFi�4B���x�RW
�u7�����}fD�7�Y�F������	�棔R�W��׭4���e�)>&�<���aG9G y�`Q�ƖQ�H;���B�"��ZQۓç�,OR�־�SB.Hy�8Y��t�U�#�[��a���NO�|��}�/WW�����o�������'2uFdAM�3��S{�/i��&&'q.��Tlmo�����n\M��J�Zu��;�B6�u�^��;H
Du��s�S⑽�$@MU5�ZrF�(	���l�<��� ����}e�/��T���m�F�x��e���3�h��칬��xhFT�e`u�Q�Rx������3�m4==j���7[�	l�G� ò5��8oϔJ+[��|�����<�2> �]]���D)�!ss�SE�2�E߾�;���V8:9i��%����><T41a!ƽ��/4�������sR;���Nm�N���߁�a�;����$�c�����Z���~��=0܄ǡ���rN*����U1}Ђ�� ��Bj�i:<��HR�O�M#��ъ9F�ddF��`3���V����{59ƧD��=�����7uw���#�b������53|�T�ם~]y�/�6�K�2.u���=�E�����9���|�Eޤ��B �zd�G���4}d��x����]��#'**�O��G�T��� ����yO�X�5ɯ_��K��u��`�J�OD`��iFF΀A��.��6�o:,]ԝ�F�ZT_qCV_��:�U=f�ɞo=�;̈́zf�)T���k�+��Q��4�Խ����&���w���I��}y83�_)G0/��Me��q��8��uͭ��`����Z�*�������X�7i�鮿~#3=�j��J���8�F�<�yڪ�LG����%��<3_��H;5���F��h
����h6g�:&�����`�ZZA�^&��$)8�Q���'�k2d���}Efn.~��F���Ν���Pf��7�����c�q�Yɻ��]���O��A9�0V���+~"m�=��JeS�2䃔���ʵ��7�4�	T��F�)9P�����`! %CN�`����8$�����9��u?A�������5����1�tD:��8.���k����Ɨ��۾�����y=�)�f��:TЈ]��}��
�`�,�N��~���N��cL�y��|[ɫ]�4I�ݥ���'��dc�/�g����k8ҹ�s?�yؼ�0��d,�XG���c��3�M��o��[�{DU��Ə�Y���/�]�h6�8rD=k��#%l�7x�D�}��Hm�gӸh��KUrR��eԡ��v��'�p���'1k[I��b�ج���:�20tI���ol͈"ox6\]B�0H+)5ŕ���
D����bXSn�{~�3_<>�j�ɡ��\U�,D$}q�������1CGǻ����u��] X1N�-+h>@�c�
�j�����Ī�St�l&?~:�z�=c⚌Å�m����y��Y%Ay�+_&��6~-c�b�����ϣ�����WX\���u�t�b�����pٟPy�.`	
����m���+{����s�`k(~Lh��Y&I�fJ��x (G�1�"�=���ذ�am�����c��S@�u�ٚ*�r���{}�Fw?e��/���?%fz%�q�{RÍ}�q\]]�n���ѕ�@��>KQ�yɉrJ��������yW9[+��ë�i�4zfp˭�����Y`�e�2��3��`��y�p�Hd@�AG�N���*�p¨!	~��.�J�wee�0��}ʗ�e��pzG���S(�bb`��@Ӗ�A)�76\�2VN����������y�z���Б8����ŕ���&C�L�t�-����\]����0�j+��4�}莵�u��N��T1ʵ�"�'O�#נ�+�kkk�	�-׻^��e��Q�8�?��U�j��:4��<Cy�lI?�ƻ��ƛa*A,"�-1ǚ$k~��~d߯FZ%Nu������K\�]��ԟ"��oq�o�!#���f����NK�E�3]��~"�E����b^:_��#F�z#.����y�~��wa����[a��U!!��J�K-zl���oݠ�/�:����f�P^U5�8����t�&��[�_�#��`��"Eĺj'd1n�d!C�̶|��c����3�Vx_��m�����"�M�PJ���k�y�*��!�;���`#�?�c	��O��~���ǀ�*�,-�̥s6g;x��ރ�����h�wa�g�Dx�����2��ҙ� �ŋ�$�1����Q ���R�U���++H������U�����K�)�����,B��s�+K�M"�H�j$4Is��j"�lk�)�@�dh�iz�w�2����I�|�ꥤ�ڗ:ҝ�����c��c`����(E	h�<��~�g�r>@g��rT�A5�'�y��^���~�L�I����<�%�\�ϗ0���R�57���
�`;ZP����c�1%�O*1�/Fy��A�@
ZpLKK[̉A*����zP���"��?vK�����[����G�h�;��H��+�-�����$o�8�����*$K�5�DC'Pa1�Ç�7P��%�	_{��&�r�g�ܷ0��/HV��!��:�~I�������r�������g�~��!a����5?����.�q�2ջ>�¨�V��D�����m�~����y�:�T�n�ޓ�U�Pנ	���G)��5S?g~AA����[O�][\\K� ���@Ǵ?C���/�Ǌ2"�q�oߚX�"����^��d>Jta�;�/#m�(�K��i� �Sw"������"`�O�����嚹�4��Z�_z#5���T�ZA��FW�l��U��������Ar�|�8���ct��~��e��gk�)��:�n���dA9� ��
?W�GG�sO�ٜs++E

�����mMAx;��ӳ۳-�Hm���S�����z��ŵ��;��W3:����9@��c����xk��r��������Ѹv�žZ�N�8Imsh�w��V�槃!��Χ�Ls{�(( ��7J�_m~t�������w:(��� �#7u%񀢢�
��V�=��S�g�'u�����8���r'���˨��-���]�Ȩ.K����g\��;����A�Q�V�;���ώw��~�B��������VQȤ�)��;b������.Y��㧇� �O_2�ޏ��ZlfHV.J�OŒ���~3��ƚ,�$���Q�#JXo���
��۴���/9���4i�,�Lf@���b닔���	��l�6��l�|�4E�k�EFF>4���.��o�ݼ,P����AZ@"u�r�7��VR=�ӀN��c31�쳮���%���y� Ɔ��VVQ)1i�Z���w�1���R��N���s�� zZf���x뫾��+L�K���\��c^�7�&��aL�4
�$ο,W��]m���x�Xx��-�B��x�@�uǯ���7��]����_{d��Ccy�W�U>�:��72�ԯ�B��!^�TO���j���9��8��@gd=&!�y���t!p��~W���q�З.�"j���W8���+}��S[a��_��.v&��x�^�k��=As	

*-�>I�_c�5>�9Y�P&����{������4,4U5���)6&��A6>Z�$�|��X��e$R�u$�;�m*�2��	ȟO����o��3M)����v���2�y��.��0<��K��L R8[7�s�w=�P�ZZB�&�� x��Z�ȺZ�Z���zx^��>�zw�ek��q��+�䘔�|��w|���85'�PR���W��������5�?X%ٜ���y�����*��>�"��٫���XuY��Ae�"*fd��6��\k9O6b�?m���!rW��#Ğŕ��o��_�R��ն�UR4j�g��{(�����88��b����>S��9��G��׽�Fڻ��|���߶�e����� �2U�ϵ9��[W	a��JD	������h�Pn^ޫ����Qs�yyy����!��!5���H-T��폽*���_|��������MWW1���!
��<�ƣq�Ν�g�`�Z��1M%�Ji�${���T|r��j��9��Id�땃�C�&�a��Tk�􁴴�2 �}�.�it�n~�����J�C�@��	T�����8h�l��I[֩�ڧ &	E�7�����	� �NGۦЁ
	�߁�rg"��dM�C�Y�|bb	ΕC��Ɓ��:�z3���L~w2�࢞���GЅ<�00ں�ad�-xު����z�B����<�]3
����=nh{����w�5��������$~�4�����[k�#"���M�Dt�ӡ"� ���Z��*m��_C��8����-���+�g��+4��1i��rt��K7�q3=��X����m_av~����{ݭك�I�S���8��;���Mk��f���m��by��^�������~����Q�'��i�4���h3T�Ԕ+�[\U�gY�7=�M�lo��������4i[ND���`��z�Ff:�:����K��8�3I5�W�}�Kt��~�^�{�OZ�
s5ş���U�$Q|�`��(�~�ao����n������4r��&|>�n���7�QhXS�o�}�!88��N7(�}V�^Ó���|��
lh��.!A�= 6�迗���]�{��Z�)sL7�$��\�62������������Y�U�S����Y��+-S֩	�i����A�g|S�/�z��ê�\��w#��1���m�H�u$&:���E&��S��뿄��Ctq�-�ۄqW�Κʴ�[S��)_��'#@�-��Dy�W�[	`�<��Y���:j��������?��(�DXu4t>M�ʿz�:Q5�����Y>��� `��0Z�����0�Q� ��(�����-0�	�X(G��H̪�Q^iGL$$���Pk��B^��:؎�Pc�y|XY�$i�~?|��}��K&��ۢ�v����=������hk�C���tb/wX��v��E�K8E�=|vvFNْ3Bd8�\�
<�(0l'ܨ�}����`H�]�;KʧN1�&��.
!��<T�y�{��P� �h��|?4�j�����h����#�U�l'�ǉ��$v�f><1����P��.,X_�Z�����"�]��jq��/�:�0|)/�i1}���6��'�c�M�@	3$W#%�,�[�|�WN%�M[���K_�	��W>v�ѿ�ee�'�da*՝i��v�gD0�����*9}b�����K͒	��nsh��lG�:wux4@/�;_#A��B�V/\�]�h�~�{��v��t�u�|�5GK��/��g#bG�������Oi��XP�D��}���lh*6��y��׽:G�J+�ʥ����P�|X�~�9�X�����fm���#I_��*��m���999A����s��R��P/��+�.eTN�W�+ڧ�;�ƺo�L�#E.�t��{AR�,�þ蟄.ܵۺ;��"�D����Z���V���JK�J�a����`���C��β#���a�.�;5��&���{����@�Q��s�ďꌽ#V dpo���ԩ ���x��Wc��"h���}�I�|��������n�3������A�����Uϟ���<�ĜB�������_��Ӽ�,&v�%�UZ���)��*so>3�$���U�eP�`�`o���9E`������F�ۖ������G`����p��" ��|�~=��_��
�DBo�PY"�,f��0�N��tCq޴�$�e�gD-�����?����q��J����?dV#�X�9��ߠ{�(�����ⓑ%�X��Ru��I4�m�8_e~���Xp�Ǖ-�(�{��(�	�|�tg,(}�'�jH��p���z��O�S@���z|c���1KH�%ũ���aa�J�y�2���}�b�(�Sf��H��������� ��n��TˋM���W��Yc����|���ry��S��Q���_�@[�3�]�>�b͈_]��qT�
y�ܯ6�z�h.��V�.��=<R���U�B2��o߾��=DMM�W����S�$4Ĩ�|Sf32w�dǀyh�ó��G�LrΜ1X���2�Y��Y��~
��<@-��oZ �SqeuwCȰyߥA4��EfƷ��)-��7��IE�Dr����r��p�S;7�ӥޣ�=Օ~�k�u��������C��HO̭FJ�ۃ?�!#�q�<��0��v�	B��!F���Z,��.ǥ�F�q��XL[.�pjȽ��3��Wc��u��.���g�� ���hllm|{٩MQ����?o%�֭8gy�����-h�U�ͽr� ���c8pz�S�����KK˙ GkS��wj�h�-�1�笡Q�ѥ	�w��Z9�����!*H�L�_7l� �|Q����q��%���'WR�`�-����=ci�4j��V&&j��N�f�ȡ�V�*��Ӽ��y��4����m}k?�k����fH�
�r��͂#�7�kCy�H�F�������t2eeez��U�"s>V�"�����(�)*�@�Q���[F�i��fB��B��Ӻ�J\;W�eת���GV�j�>8m*��~#K�A���>C4��J��SA��]v��g�<&T`����@4�����H�x+J52�ii����o\	wh����N�κ�'�a�S\�R�uOu
Q[�E���U�U�:�n�a�2��|�8�:��?�t��D����Ƣ2����,*���Ɔ�Є�̘\�v��VX�H��d��m�`����^���e^z�Ե�p�j/H��ǪY�m`j{9���jYY��G�W"��޿���-Z��5f� �0��Td��; ��;�Ξv|��&I/��b���㣳�����T���Y��=�qߤ紁*	Jf	��8Τ��儘{ҷ`���l��>o(�o`do�>5��j�M�{��K<AH��������2�ӧ8�>�*hR]��a�������	��Z�������.113+����1�eI333�
�����C\��ݟ�	)((��1`��A���j����q���
�T�<��Pd�mߞ4�+�6�x���г�ӗ��7/N-��Ð��P9߯�f������5�㇞H��OP�����5�b�c<��]Jr0.=�E��mYt��,W����)+7^�� �#oz�@th�
A���Xo�(�2�N|�U�  ��$x�懡Эɰk]I�1Rנ�����(�d]_�����;�5X�14�[\� ��S@��pK�յ�����B�0I�U8���`�u����~{{�?#��yb���KШ����ݹ���*�����T��ڍ�e��)�N���hmm���Ȉ�!sۚ"����z�$t��2�}W_}�� =��_o�"V��ĺ�]X}��%kB�Eæi)x���f
Yq�H�g�h�ּw'�*�V:�����W|����߭��:���(�U�:c��ܴ�l%�@��O%�7�H��l�s�Tc�/��Yg��g�Z���炌L�] Ș(a�%8�4���<[�� �H����n/ǘ~9������������ܜ��X����ˇ-��7B�df�'r+����L2�e�����_Ŝ� �"!������~�@-��>�1���ɐ�����������uMgaiI��{r���5�w@�0�C��uS������?~<3?���3tk�0�����+Jʘ��R0������Xu�BO������TV�S��	�f��P����5}?�m
��QuUֶ�р		;�	�O�=��:�[D��+�탶��<���|�Ǵl���Ry =�C���^��3m�:G��$��@Y���Rk
�6&|Ym�4�j����P.#��i��jO�����K\$�N17z+��;)����T�ޅ��Z~�K���ᣔ:l##�=%�y���@N�Q��/��|O��y�6�(^�,n��APX߽{��ty�N�eY�s�ã���Ƥ{f��Ʉd1�C�F�`��1|��XO�>��ݵ,�!e��R�w����<pHOvO��l��]��[�@>$v���������-L�u��կ������f�M�/O�R��0� �T�@LD^vDS��K�a�m�od�F�t����4?Zz$�m�U�8�0����G�U�ׯjy�s�L�j1�k֍�o��G���q#4Oʖ'����G�E�=��p�2H���-?���Z�L�~�ז>���̳";(\��O���"��L�^hi��0�xˑ���
&�I�% ��*��T�/��Ķؤ$�ɨ�����iy���-��A���3���?~�7n� �>�1H�LH����K��_Dn���2��k��TpUTnе6��}�M6OS@SYsJ�_;��|�E�^{>���͆�����E*5N^�t �wwX��p�3hS�Q��9 �/��n?6�҅Ylv��N�5�G�uW>Ҋ���B+��[�����|�9I�);�r�-bq�5w�T���_{�Q�����;�&έU5�����x{@�f�Οvly�T��S��ĻE몕!�b�j#�D ��'f��TLL�����(��2Z�TQVT? Q�['�[�^_�	����s^P
~�:�����*����-@�,��:��I�RC��c�+��캶AJ�.	i�.鮡T@D�)Ii%�a��R��;���A���?7O|�����d-\é}���u�s�3D.)�t�ʷ����5;�(I���OF��z��%�������<��s��b�HƙR��W�o��1���9��'��8���P�F�&&���`7�M���h��Y��j��F����衖︍&�/���ǥ�����y�x�-g�Ҋ�ޓ�FF?������0~��0:���D'�]����@w�uLs�!��z4P�Z�tm����5ϧ@�����;C����?s���
�3[ZZ*�T�����=2ؖ��Ҋ@���*�-MT���ݣ�������-M���d�r�p��|�%>�^�u:]>�t�FKs�,zW���	7�h�l,B��;�8�9'���PC���1�3o�,C����󽎀fT�c�ЩO7��Չ�a�΂���i��!�|ɰSu����9��v�o��q9��U?�Ed�D����cX�ϳ��X��#���ȯ2|j�{�VI`���f�z���R�F��"<h�>���lEz�g��ذRRR�F$�wO�q?�l�~)-���Qu\�:��P��3^�����m�����4����ZO?@�݅o(%�Ջ3��\"h��H��~�괫p�����ZM�X}%��/��\x� &-w��S��){rM�W�1����������Z������sx^�D����u�v�?!�v�!�W����p �w4�cA���~���h9ٝ8��ԃ�����q�[�i*m�͆�����:�xӫ�7�u�����G}Q�{��c��O����Ĉ�Ӄ⃂���w��Ξ6p+��+m��՛B���O���z�J\�6M�G
4��X���kn���"S�&1�9H����?عI�ft�0���Ɔ#`5��dJ��r�����Z)	����3/���������44H�h߰j���Q�|�7޳�Ҽ.���k�n��������ۭm�3"��v���_�a�/r�ѷ����<b�H.h�N�2��DUͷ9�B����@87�I:a���d�b�>2�}:q8s�Ւg�_[���RI3{� �f�sI2OzĦϺ��	3[-qw6=I�T�`@@SU�#��NdoH���G��9�n���{̝�0Xc>9�T�4xcqpn��||�܆�zv����	=��[Њ,��;�� ..���
^��TQE�7((�J[q�?��!������o�IF����Q��mYߠ[�����'2�������OJMݵ��{��5m�{���|<i���t�9��_������i�H��$;{$9aюl%��v>����"��}�	O����f�g�߮q�X�k۶��ck�'O��w{$�2ǭ$��}[G����ڥin&���x\�~��I�t��9�`<��כ9����#Tt剴�l>�,j��9=����Iӯ���1��sf�M֫�4�6��{:�o�5���9·�rs�����o��zE��AA�(��]v��3/��sto}������x9֛�@8VN{�l�R���6}�3����a7Q�����WOܵ�ʺiT8��l�v���ʟ	��̓���8ը�Q�_��J"�INƕ��!.�G����]�+�y��o�}����b�(-g�������g#m?�dv��AfG�je�a��������c�Vt:��ʮ�CݘN1��5s�n}��2{�|���;�眮h����ͦ�� ,�Dߘ���ҍ��o�گ��dVX�ڛ�.�ѷ��d�@[����v�Z�nfaR������4�S�99evc�}��l��-��rrOܯ�ű��H�??jeeu�A'��4P0]�̕	�T5i�kWv���&��Yt�ft�0N���w|���&��
�P7��T���yO�u�F@<$���������4�K�C��6m t����)���{��'��ħ�qBc��빯��G���f�4&+�.JL�PZ�ܽw����=+���A�uoѮuӁ����i^nN�����B���0s�-�ev�(\��X���t􉾁l��T���9��a��7�]S��׷�2��FϽ�v�Z����\��C�B�	����uY��=��k��/�^��J�Q#ф��g�^�L�4��]0U�۱�Ap���)�]��*�����*O����n(k�:�E/G�K�1�v�ew�!�����u�-��˙��
�����8����dH�GW0���|F�χ�����QU���f�;e?�b�9����"��z89�^�kt���\�y'�Ī��aa��Z�pۨ���ZxD0���& M���?���8�Ag�;ts��rqc^�8}�v�����?3O3f�]~CM�IЄ̈��/�=�8��{l�!0Y��EJ�x��r��	=4�73=i��G����B��;��Ѵe����C�}<����޻��t?l��PSu"��n����V1$�S)k���=���G���{����hs�>�0�χ��2{�o��w2���6a�|5��Ľ�(��{�SqH��H� �%����U��~ɔg����:>9)��x�BRw7>���x��X�VʃxvL**����Qk+����`ʽݞ���~j�s<�Y��]\i��dOiA9��[�c�b��fsy��׭���fL�%�C�]mY�q�m��Q��k;�-(>�����ɈSɨ�5��n��(��ʶ,Z��ڽQ\���/�	[���߲pcj� �(�h�?B��)(�����20#41W�E�K���B��py,��6.���P�t�H�=v|�M�sM�P���T�D8c���1�7�Ǝ<�T�Rr��`�Y\�	$��q ��	���}�Ŕ���y��Sĉ�w�8=�%��[��gL{�o��'�����&��!����̇.|���8�c������H�����4�{�\]]��yQ��J�z����--O�?�5= :�sq;�^ҳ������?2]�Ԍ�C�UV�����J:u҃�ڦ}�6��� ��+W�U���m^���y.�=��=����H*��6p,R��Y �У��Iߴ\��Jj%���v��/П�&GZl�U _�|���S�c�C�ӕ����O7����q�tE�1��
*a�O��c��<؈X"�+ҳ*��J���I�ɴn���m���Ht����(��'�N��Y*�0�5������>�C���B8N�E���@�~[�§ ��RPP@��l����	bV�ٲ�9�=���"�1��^�L0��q
�F��^b��:�(j,&�ԛD���R�A��l9��퍤{�F������`yY/���Ni��(nMU�Y:��5L
���w8��(5_�j~w�q���h��p�6D�8�a+�&q;cH���)�3�� ���Ha+�����K��Ԏ�P4?Vг\	��Rw����%k=gs^Tkb��ϥ��^� x�Qf�Ǳ���FæWB�������q:��V��i0��qԬ�F��)(���\!0-"&����J�����:	�Xw���y���}�c%_�� ����M����)ǰ�eN9]׎L��+�V�~F�0��,���W��~G�|[��ɗ�r��G��1N07x'\r�:��1���-q�YCS ������.B�ӷS ��B�ÞEsݢݮ,UV[V$�L5���F­�(�5��R�.A_ `�9S�v9v�WZ��,*G�} �28�zh�L�����}7���4�x�c���5뼽��b���W(����
q@���� �(�T3ߺ8t�����O�doZ �C%���HA�#�B�vVx���ٍ�F�=��RI|F��wnJYM�<�.ծ�N 3�䓲0���miad�>��b^���^��g��<R�'�z�¡I�}!�'���B񎾿L���?��D�.Ui�yٖ���w�Q�|����aVZM�C�k��3����6?@`}�c�ӯ��4�3Jx�:�|����߭�%��j�K������lp��G��޳Ñ�ΰ��X:<��&"P�E��6�`�x��̚�֥ͪ��p�pޫ����;�sʟ?����E��nZ��&"9)���s�V:ך��gR�V� ����SD�u����2و�(3�IǳJ��u3+;�x�S��ϟ,���Kr@����z�_�Ƃ32A~FhѾ�qT��ф���w�Tю�������:N����"s����}�.#�.G�X�SI��hA�$�3���-� ԃ�k���r٠o��cA�-�9����tv�LY�,�Zv-�}��4to�b�ܐ�����Y+��e-߀A�̩D8�����O�ωOQ5Ǖe���%��!���U�E!w~�1 �u:0��%���`A�wO��Y>��u��O�OW>(�(K5�/�/z�N��!Be�|�t��h,���:3�}��f뇎�5�8^G
f{{6n��� �-,�b�� ���g����Z��/^��D� �K��Ug��T���j���CL�H��c��m�~��T��;�S�5M �x�K�E��[�3GWI�����3�oi�]k�����(��K�)��}�+�}Uo��ܽ)0IX�Ǡ�q|w&{/֋���G����c�ښ=��&V�0�)��m��0tά��ߣo�>�A$(A�T$
�Cы����x��M4������$���]�:^��̈́)=�*Bf���2�	���� hv�?�2X(����)�|��_Wz�=����cI	5R��
��0@�w���]a��<���=�<H�a��s��zo�۲м���+��NL? ���n^��]�	�Bk�� ��c�~���gG�H��F-K��p��Zم:����N<q�/@sNŜ,��Zf��z>���?��KY��ڷc�}�6=}�$�F&�d+��V1���,����U5a��I�����B�/5�0�*2��������uc�U�{�[e�^Ă�}5�e�|�L��FN_��2&XlF�t��u������>���*�}�'@�Gٲ	+�9Y�]%nȓ2(�>���؈|n��pp��Ѹٱy\�̌���x�D.
!l=��mk��]��Gj䢲���L�('/y�����y;��	Q\*6��M���t[ �O�t�z3$C��H�d�p���_!��ll�6��I1V-$"���s���0��e׋r���%��0�z�ذ�G��-x(@	�W�αJ^��O���n
lF��n`�<.�E $�^���-l�]���y6��[}d2ez�j2}�\�\�s�
Ec���;����W�4%��_����b��&���G?�k45'�j^��D�����g���V���R���ϗ!u��/���.a�,�WM8��.�	[�0	^��R�>je��z��T���I���bqq1���|����:)�%h�.����xz����ެ�P�:R#����]]��Xd8l����i[X��jZ����FRYl ����H���qh��s�4�ʡxb��xba���u�;J��Ⱦ�m��G�_!�"]qc�KN��E��{#1���#E�o(�.�n��3����yY����%�R�)"fV��۟S|��>��Қk�^<�R����υ܌\=��X�K���$��(���ˌ]�F���|j��Sb?��ݎ�أl=��Μ�o��5ۑ�fEJ�9������ܲ&��4 �� ��llHAȃ���Ζ7K|���nei	x�cKKv��%���8�{j�]���Ҍ`�i����I$�?��t1�V���>���T�6_��ݜ�����۳�k.��0� ��ƭ�	���Q�������|�z�[�cE.��Є}5U{��N���)�!�~}:�����nq\R]#�����e��S)������a����-1���p�y�
a�R�r���;,��|U3l r�9���*�O�Ý�~ݛnb�Iz���z���e/�sz��%�-���j6,�w�u���!ֆ��fE���"��A���`:����',��!�εX��*y���7}�<vE��S���8L@5�Ʃ�9�����%˞p�4�,;z�y�8�v��t��
�����H��֦����x"�Ŀ�Z��%/�����ss:��l�v��_ۚ��a��d�����e*DƸUJ�W7���.������[�����P���˫nپ����ܳZl I�~��-�ϲ���~�Y9��3Hs���	��'i�����;4�ӻ�2�ڄ<z��{bZTpii�u�&�b�\� ����kՀ2�S%�����E3��%�А �NAA���Mߊu�#���%w�0k@�>���p���Iq!f^į4�ù����]~�xu��ub�@|��k�E�W�hÿ�Fv�җ]8�uZ��?���4s(�.0�-X$��Vo�}�H�^Z-턘�����o�?e���;ψ�B�+2L%�6��{��|~�ӶMX ��S�6w��5I2+����L���5O��S�g���gt��9����>��r�Q���c�ҙz��?�X\���v/-N�Vʞ[K'q�,�R/|Q[}�[ɧ	UJ���Z~����66>���>�H����噰�A���u�����z*$u<g/�a����9U��ڶ�[��3��4�Kj��!�r$�e�� �de�I�3�~.�;ZCCVK��`ʖ`�4:`7��~^��Ҁ:�W��Խ����){�JR���S�������0�K�z�ėr
�+�p���Rp�8ѿ�ym���&���O�7�I��^�h�V�������&��}��?<��:<����8�Ժ=�����gwJ� ���[�^Vx�,�������?-	�,ŇZK���}�Qh:(Dc/���n��8"��5�;��5N0".�U�#?TWSyyy�l)BGu�A�S6���ԋj���-����/J>��W�PMP�w��4���
w����!�7!a��EL<;���]��O�G���M��D�-��dFOci�p#�7�t~'>-�3��iW����c�'��H�R���t���M�a��W┐�I� *���VU�q)l恚�V���/�:�N��y�S{R���}&��#90�E%����Ԉ_޵7e�.%&)ġ�R1����t\+�^&Y��Q����M����6�m��)e����CK�4�I:�~p5�Pt���w�æz��)���%����*�ҧ��d���1�k��u�c�{p�ڌ�H��&�׀�����*T��d�T��ƥRrI9)�а��S���a+'�P�C=��*�w���m��3��
ӡa~�.��}�H-H������������nSw��k��3,z�B�7��k�Vq��:�t�H4;m,��0���MJ����uy��O�q�H�����1kuX��x�70okt�,�ǧ���ʖ���ͥ<pVR?��~{��pw�(L����ăɲZ˝2޷��w'���T��9R�?*D-�ϰ��c����]"|g�A̭��I��Q�/�	d�A�:���ul.���\/�)y5v8;4�����_�\���;1d�C�m&�I٣��Q�F[�+����."�<����?�a�d�U���I塜ݱ�N�oR�s�O&]��%�E��j��k�(F3�M���mL?�O�^ܑm�u��:�b׌�}���k��R�%J <����KŴ5�,�Χ��HǞ���U�Ũk�򻛻��\����9پW`�E\�)�1�uNk-3~x���|�����	���0��}g`�-τfM�[��&�լ�F�-/���	���/��DE�o��WKlw�t����TU�E;>��a�NսC��Č����^a]�,�es[���:������5{�!۬�}��L4� �(���́��#;���ΌJ��'�B�ڭ��d�|�( >![�o���!��5M��ׅL�
3� P/z�bnA
$���I�p	wn	W��y��@9V�K�-�d��k�B'.55�QMkJ-ʙJ�L�uf�(�k5�A����)���ӭ�t���Ũ��h2d�'H���1�T
�^���)��3~(J@�22��`�h���������,��k��I6׽ﳙ;�%���z<�r��F��{r��P�#��7+m�>��$�|R6�܄D<k���bvO��e�Tt��2l{Ε_H����v?"�H������bg:ɣF����(wW<��]6����ZJ2^7�TzmZcbp���K�c^�y��1G�m�Wt�^�]�yߐx�J���/���h�����)��� �my�b���?c弡,i
.�@�����"�G�#I�e�:�y���A���r��!�����O�7$�#��H�L��������Ԑ�9���+�@TM�/��Ě
Gd��k�Vr,�w�%��V�Z���G�RH46kΖ�E>�=�V�i��+]���Ӂ�ܲp��_#_�M"$���*��T	+F,y��p�veoi��#BnY�h?.��!�K�g��i��QUs�SQs-�����l��T~�W�Q�|���u�,=���0}$A�m�52i{��5W�C3p2ᾢ{36_鏘����{~�L�;r#�DC�U+ӷS�K^ߐ��\��x2�����l}��+���G܇��"J��l�b��e�������<�|1��<�E��T�r�+/YM�Ƒ�
�kF�]��0@Μq�8u��K��Gܞs��E��S�	������5m��*ߓ z�����J~uv�7MD�7<�*�* �!RZh[�z}�$�}J{�N�G�����JĞ;ȏ�!��R�~� BQ�����=F���{D��]�:������L�i��鼛�Tq1[��#ED�L�;?{����^���v���<��onKS�FʥG̾UujO7z��Ҕ�l�v��x�'��=��io*:;�X�X ��w�%�)5_͗�������u�$\�-��[4�"�h�A�\8�r�����whep��ܷ@�T�������}1EM
�V;"�#_?)��K�������*�(��'D����r�#���u$�W�ݬ���xS{)����mv��w8L������H��cg�YGN���qG]g��	
H�uA���@>&$��N��
��uJ$e?c���p ȮO��+x�̈́ٸ���a�o�I��uӐQ<�j(���]����FGk��utJø߹I���J��!B��6���թq��(Uu?=>��y�Åm��)Q�jq�Io�ב���o'�#*r� ��3�W���qun���&�6�G�A"5�9?vҩ>�:��v�	Ju�yd2�����3h�юV�C9��t'��[��ʦ/������9MXˉ����=Bn��د�}�c��7hP(�e0`���#�� rs<�|@==:u~9��#[:$/u}�T���h��>)�H;���+&�Z�S5>\���u`��'�։������sxz<"z0�tJZ�fm7+���"��9,�̾��O���/�"�"� ��V���Yg����Y��]<-B	��I�w[m�����4�6eY�~����A�w���ԍۀ��=�v��p�����B�v���
��a�A�CE�P���V_9S��EB��E:�!�,���s�4�E�>] U��tD�2S`Aq�(@�W Ջ�P�|��%�|(�]�OW(_ݐ��+�z}����Ӻ	�8�v�����_���b�W�>���;F}����'I�:�?�VR~smO����>� 0���Ǔ�MI4�5��s�H�����q�0�]�J>+���~y�|��k��/���'Q�V|���R���߻���c�(#����A���j�ܐ`H�[�������鱌2�%Qΐ0v�|ޅ���	}�w�I:Dt̕�S�LǾw�%$
��E�e\g{@����ɦ�G�In�q3d�z�)�e�H��4���p�-֜�g�=�Ҍ��#,Ι}ݺԡp-��L	7"���ܱ�1��f�z��$�y�T���٥+�}O��aa��Ӆ��`H� �C�z<���ʅ�u���N�]�~WMf�l6�Y��[G��-�����Ƶ.�!��������di��^Ak�m��~�hf��:Yr6C������a�����_��c�a�@���C�B���2���F`_���{�~�4[�Lf:a0���Z(��d��fωMɸb�Y$A_9\Ti�4<��D7rN���MqIq9x6��z�9<��^�+�j>�:�R}H�^qb�(+�ݾ��O$����bO�s��^H ���tW�)�z���4�p� �?�:	����Bc�38?>^�Cpw+���j�þG�v��pH�qڨ�R��Q�3���n��8v�0���>�����_�ޅ��AVI�I�v3��W�:�A8��hWZ�z@�{�
̮��J�8��F�Z� 4��UywZ(b$�ާ��=�st�<��}m/\��o��xv�������>���#8�n�K�T�kY|tㇵ)�z�%-���;��W�畞�O~�#C�(o����Xl�Lc���;*@���_D�ʕ890���f%�� ��	��ٗ�ެW.Y�gƂ�������5�5ȯ�x�#����@���������y�׸8�A���6>y"�M���s�`j.��}U�<3db�0��T������$&y�/a����;y��E֓���r�K�Jf��aX���x���aJ��J1=���lc�l�Ӄ�s��+����άC��t�V�)��6��^������R�w�G�G5$��-��%�<{��L(ɚ:�1+٨��7Jn/�ۏ_�EO��Em�ʢ�6���>��9��(��pg���j~;���Q=�_|n���6�&�N��@P1�È���0v�lcT�Co zAL+GH��@{�X�B9�	�߾�vT�HV^��8�+y_	:T�e�b?����iP�Р\]LJ\�8���w��*E���w$ɗ2��&hMԔ�M����`���`Z	��j���տ%�.$Q�qW���̺��i���~�4ZˌK��m��W����B7�R��������<?<��X��֮Y,��z���DTl�2�|B�Q�h�P=�H�w|����7`� =�ܾ"HO���S���2|��~��ҷ�I�w@s��T�nNn��"����|wV'ȶxZPc�|����IpJ�B��0��~����Z����`׀h��7aJ�E���ޖ%�"_��!ucQ��d��L���pr��
`���Ԩ�0-.���%j-h��i��ʺ��k���WFo�L�LW5O�M҉m�/�3�T(��a�>��h�ف�Ehe��,a(0��z�携o�z��K���#�eP����o��S@PB�ʎ��)\%�>�		�(e��	�gKu�S�Tݧ��5x��(����7w�gYr�k7��`�$�-6��j4%7��M�ě��G�r�0���h�_�\��($$��*ʮ:��giǥP�L�S��=j����;ymk$�78�⟜�8	'���Et����<����zR���M�`�Ě��NŚ�D�z0��Q-�e���_#{���Ʋ����G޿�M Z�ޭ~ 5U��Xl$i�h��(v�ss)t�l4�N$����Ƀz�Y���3>��,j�n"�{��9ݝ'?�<PV�I�3��j5t�˔�����3��TLj3��;���T��b��������a4ߥ*�ޱW��fP�k��%��q�2x��?&%����
���u� t� k���\�Zx�iil�
rۈСh-@Y�>��B�O	����!A�����y�<$j�:���p��zV �}93��vH|�����$��_�t�[�� Uo��g�-O��T�ri {!���A^���9�D��C1�s�a�`'��*٠;�ldW��0M����,�}��Ǵ��+�p+y��O�,ioW�����fx@�I�}bt3���V����8l�W�eϠ�O��>n�Bt�@E�S?�fj��y�ة�+}Ι2��"�!4�囙��b�S���j�t�qj�y�I'QY�v�⮸�%S,��;P#X`���w|� F�tG��'��6w�륻�j�&R���ɚ Dp��
]�r�+Ԛ�p7;��̫�ꟕ�Dj�P���Ϧ��z|drd��A���=�O�p`���s��D}�^�=Qx<��A5_=R7t��qm|gI�s����d�$_S��B�S*%��B��>�k��g��~F�Հ�~&����`�H̋����v;�̴:��5��,"� @��pD�0� V��_X�#E��)8�h3�#�pW�P�2�X�^�p_ma���~b@�-�I��F�bA$���ֻ��/����7A?]ې��|���Qq@C��q��Z]������go�o�mV��䀹U+��9����q.��.$ CC&y����-pC�JU:��M�x��F��\��D �'+����!�s�K�6�l���l^n��2�<���^�_�I��d2D!�`��z{�&�z.ʊ������!��ˇ���]�c0�f3�s^*�N�B�qE����h�̊���	JǋtO����h��NeE�t��T������"IY��2�P"B�[�Ow��r�v��2�"�����??q���s?.1��M+yiڬ����uEz<Ж͐_�w\\ м�	622��ی�<��=~���hS�-&��V�H�T�ID|3�k���gO+^M�p�w� �tn2(M�7�H�c�9�A��1���Plb��b�q�!��w��j$�~o8~PXK1����C���my�`T�&Wြ�'kM2`h���Հ,��� ��\8�IT������X�z��u�H�[nK����I9�s����x�R�\��wX�㎱�]V̩�g�r�B�	����PK�#�^��YE+S�w)����JNtfTߨ0������i���a"zӆ~�9��QǝQ��� �7}��A��2%J(�c

b�N\�6��0@����6�����L�XlC�؁X�z)(*_:
Ln(u�v� y�.�r�l�I�
���_��� ��5�B�k�	������/��"IW��аTj8���B0u��&�Թ���^l����^v:��A��)�f�L:^���;�	�7�F,VO�x�*�u�ޕ/x?~���[��8���3tB)a�e:m>N��m,�$� ���&�q��U�� ��fv{�]2����lQ�KA�����^	�^��������F��<�G����\�z���WI��n�U+u:�ª,^:��ן�x�~�DI���� �3'�ȕbh����1��uV�ꫨ*2�.	X��K���tw��sZ
,
�X���W�y���H�Ǣ���&��"��n���x2�.�����M��a�����Ah��{Q&>�#���=a���q���Avᾄa��*����H��A�ֻ~�B���N1{.�	��"r�
D���vd4���N������v7���,��<�PmO\д.gI�]0�$c}C ����ɋy��yw)�H.nn�j�'��A���s.�tC�"]:k�r{���ӽ��F�	��֥���F+o�¬ÂE����9��� My���@Ǭ�3��\Yd/T���� �..#��u����}t��)&pP�x��[�[X	й���E�q�l@qaaK٩i�q)j�q�����irG1R��b}����Q�6R2)��+�
ʩ�/^�p��_����Ύ�����`�y9t�C��
Y�+@M�����v�J�vk2B� ��(K��/9�IX4�F��)��{�봈{�DH���P���8��)�}���"e�=������1�ӄ�"�/]����>d��{�E�{�-���!���7u��sm���c���]祐�Wq&pc"ҾD���Mͷ���UY�)E���0+�����p�&''g��a����GcC$e��%�x�����>c��Rc��@7<7��m�C����8)�E��R)F��^�M�i�֏(���4;M�U� s�%�8�`�;�F�D�a�ʵ�k�?�}�A���4��Z�p/B*��_D�J{��D��kӏ�䧛sm:+`p��1���e���
Ea=�4ȫo���V�W�Q� �2���ep����Lz�lt����P�U
�Cq���Jh�����ާS�m=������!�6j��Ar� �"3m�&��L�v�b.��Ez���Tu�:�����׹a�ʈ�:��(��I47��a�yi��ì��Q�Z|�G���Y
���kW�|�F�*�P�h�go{{��ox���i[�HD7n�W2��D)�b�
��rt� �G�M�Pa��[��wN�Bg�83����#WQ\����,�LM3є�����M��c�v�����|��6b �6�X�X[=�*g8z��Ά7����� �1���X""i[a�����4�J5��W�g����x@��+��f��aD:�}H��]={%j�J�$������;��2���ip��Hп�`M���}�x��Q��蟧��+͖�J�	��me@ ��:�.ht���	�9�	�.�.�Q��/�7�^uӚ�պ-�.����G�o�Z�Z���3&'i%�c�\��`J�&J�q�W6U��ɪ%����Թ���p���!m�� {��m�4&3��`:RQ�ǱV94l��m�r t�D�ldѸ�S��Su��i���?i�_�ZF[�׷�Ps3��}�
g&D�M��^��|z�f$���?QBW-��$y�~��%v_&���R÷*�`)[^!��{v��'�:!ۂ/0�0h�I��7'����M��ֲà8�������Z�xK�GvH��s�K\���.$g``P�ԤB
�$$P׍Zݽ{ȗ�1�NM�_��k�D��dv�x�����Fw���><T@r�w��
&P��霻CSR��d-��1��"yq���
D�kᎤ0~ݬ|%Lnh��7���dCk�3}�pj���z�����y��
)��8C�����&Į���E��~�yF��Õ`_������8ǫ���U������@��ih@�����;����}:.M�i}}=G���z>%:�q����ɱ������w��	{'���sg�9�=T���i=Q",H�Ю.����֖�piHa��!�����d�(-�+P�����I�xN�gW�F8/��X�zR��k�|Q##�+�A��"�J`#��_���#�׃D&�������[h<	�4˔7	>���������QB+;�v+.W2�F��Ϡ."""h���� �[.ήe�&%Q��<��PQ����w�.�]�}''��㿞h>7y�k4V����"��?����^)���G	-4Ao��䏲�^�WR�bna�b}E.����Q��R���~��)>)�Y>��c;� ���xw�#'".qy���y`Cؘlgo�:�����V4��A,��ob(�7#�À�\~���y�ɠ!Z|���)h[i=�����Y���W��?�|O���6�zc�p*��f��9���R�����o~�A�^����]�X\B�VRR�̰f�R�xH"�ul���S����V�y���M)�K���`��X�������H!��]��.��w�F���̀���޼�⎋OJA8=m:,&"t�&9쿟p�Hh�p��
��8���$0�h�5��#"X4��	�EEAC+�׿���'
�8S�%Z��8�`�Ä�����ݫБ��$Ѥ���˩������e�Z������~h�͗4qm�����3^�3{�V.���f��^��%�I��َ�t#>�Y|l��Ի�t���׭瓼�'��<K��L���Oњtx~덂��:!�/�������V^o�4K66c�d��~���-n�o����r�~�M'%%���߅�b��XF�1Ա��߅w�ͼ>Y��EWY߇QQQ�L�x�|�:n�����D[!����7�=��#B�`v]V���o��	T\׊k{�\�O�xpٚo����A�[���<8)�{�l�h�lG�w����P$��/c.���ZeM�mc�1��V|��ߒ�W<��d<���G3��F\��t��N6{lb�7��4����~��M>��LZ	�JO�_�-���^�͗��:>��k�0��If��%z8���I�?���@;�����4)�[TQq{�q��F���.MП?���_D2�J�s=��Ƥ�oa�{uXX#33'���G��TӪ�S��ϟ��\덧_�َ���7N\�Q322����Q�6���?�qC+�.��<[̀o��v��1��[���%ݞM�L��f�[#�����R���,r?�p|x��P�8�������n�	�7������K�����-�|E�=�up������6�6�|֍���M�s5EC�tG�>�LMa�Sp� X�pdl�����xO�z��'��˶���\��[|�x*�׹]���@���^��q�[9[Cc#�gNa��H�F��R�h\�H�l���դ.n������R{��]5ϧ��?�����4��@@Um��׸N4[<D�c��?��iV`��2Dz�4Sn�d�����~�0��ZȻ~�3�/)��=n�˶�'e!���9`;�ޕ,da�>Y-d�9�*?RLl�g����\�{w�|�
#��_ZЦ7�)&W-�,�������Ao�ͻ#�s@J���{���. ��UZk�����a�}���]�9��fg}��]a�o��9Q�� e?=^OO����@̣B=�L����v����2�)����%��+�q�Q��&\5��P&�|j����'[m.`�˾�M�f�'�֧j�2dR�	���$P����D[[P��7�ige0�U+	A��ׯ]�4=�3���lqi����������sv�嶶ʯs�q��D��}�c4�')Y����[HuCCC��,|q�)������릑��me7�����ǩK��ܙ�ii��=�)��s�� ����
�
K���@�WǻU+��@�A�|��>if�;N�<�����T~��^ȋ�y�I�Зe�W���⫝&�����Ew�Hƿ1�љA?�ߵ�s�y~�9�/�g�Ew8U������Vw&�n�v�l6����ߑr�$(}v����������[��n�x��� ���:U���nH���K���ե�y\��Sj-��l�t4�t��'��,����)��I�~/��������fY�M)���AFV�vz�=�&��N|G�`�o���=��l�>eȰz�����P�S3�3���s�O �T� Jɝ]M���&�X��X��<1���bO��_���z��M���c�+O���9�ק���T��ku�H�_i��\��bhh��qqn.[ƫ���M���c�v���|��j�'��F3�`�OMѯ�G�����W����V L[[{Rw>�� �s�~%��Zt��߿�?@<V�� ��E���;ou��w�nmBB�B��dm!e/���%ٳ���N��Qdٍe�2f��Ԍ}c���>S�u����9�9�y��9��\��z�_������md��h��:� �E��^ա����/.�!�!���3�A�ف8�p�:i����lomZ6ň�	X�������7-���)��$.�:v��9z���@���Md�|��dd2�趻AY$ '���#`Q�����H�HHL$Lg���(��7\���;UH@�_bs�) ��J�Y�o�~��D���K'e��9\����
�Z�������;�w-.�����/���^�k��u�Vb��C�%|���b���Ì�k�AN���JOp�l��t�Z y1�j6�
B5xR���a��F���&�-�NBB�A0%4<<�$S���"y������������Hf]U{{����J��׭{w9���R9�� ��!��5r�s�����)�q����\�
.�r())�V:uq1�Ʃz��+ܛ���i��'�՟���Bv��-�ZZ^���|v�]�����������?��Q�-�_� "����$��=`�IcQ���nH�ڞX�$O��`�Dr���@���+�Ỳ�mu�Z��� ݮ�i��AL�cQ���4�u��rJ��q�5(�߁9�
���xLmD�{uO�ٴ&�������o��Ehá9���eȌ�)m80$*i�ML&��(��;6��
���H/|ОZ?�j����$��!��<	(x�o4�{�'@�O=ĥ�V�{�p!��{����8�U�����J��e{��K�������@��K� ak�H�&j~/����o������n6�rO8U���J\�ʥ�H7K�* '����]	]XX�"ձZ��|]�[d�/_�<Uq��ѱ$�;;�?�MO0%���1,�HX@��+v���T�E� $����AX����NK�Z$+������C1���*$1GIZj?�`�-�7���IK��/_ު�r�JQV���w�[F��\�G�P�m����q���	��!���⎄�s������@�睙��&q4�����ÿ�{̨������ $f
}7׼j9F�@
�_�Mt��ý���'2��%���- �d��8ށ�Ds<3$smk�hjj�W��Vd^���J����Ar���,d )�6�D�,�^ɱx��� ���� 6���.P^,��������lI��lu������PB��~�H��k�pK?�W~G]kZa��xKH(̗�B�]�,��^@�7�~z�����ђ�Һ���u""�A���Z������7�^ѳ�2 ���Q$^�-��4^����柡�vn��K�}�	P�G�u���]����?�?Q��� �����?�i����=�:������Zɋ��T��M��}�}�ξ�u����+��8� Jκ���I�.�N���ځ����c�bΌu3�SJ�_���d!+a��������8��Ͱ��?6���'���mn^^X�m�ۿW��~�b"+��(��|�ĵ��z�۫r~T�?�"ۥݰ+ՠ�S��S��^	0�����X��xS'�"��r��߻��\H�Ǌv��w������7��5�>f�7�	�LX�OW���3���Ԝ/FWis}ȹ���B'{���<��ia�F���Aq.����s�Zp�v3v��d�p�^"����k�y�L�ut��I���V�(}�c?��IG�U�Km�;�ַ��_J�~� ��ȱG8�i�r]x43+�oS>++�G�7O�n�BD�]����#��M/Po��F]�<��`�P7i��!vk�1"+�޳q�dϫC<H،8f^ű��e�����M�Փ�z�,��4YX�U9'�]�6v8��Ү�r��ҜL�N�;�J;�_yyЭW+���%=����J8]�t�c^��x��>��_D�?ےrIǧV�3�r��@WS~M�&�D�V��F^��@���%o�G�f�p�(�6��o��>J��:�ٺ�mR��K���G�^���=:��#rS]u�B�fQW�O}l.�f6F�ȫ�*�{����]2��V�:W#s����9�H�.�1<IH�<����#����W����,V_��=2��[{�������nt��N���ȭ���t��C7r(Q� ]�Շ%&S"�h��K���2�%��P���M�	1Y���/��#l'bq#�<��eE&���c�V^no��*�190�aD�辰�o��	V�;�ؑ�)���!���|��1ޞ!9e�G��X�v�hIA�U�B�j�׃���]�q��Ѝ�8�2^���� Ka�ۡ�B��֑�ٙb����Ɓ��m��V��+�/P�f�,E�ڇS�){ߺ�%��#�g�t;A�0���~t&Qv#�\�2CQy+�6iv�����@{����|� �z���j��^{�3��88�)����a��iᤗ��*+�y���9ƶ��3Tu�Orw%��{��#��t�}�{�R%H�Nl�%\�Ԫɭ��Y�c���3rxY�X�ꊼ=
�G��$�����8a�HхK� c�;y#�11t�u�����#��pmS��D�{~^����G�m�������Ǆ0�!�Fn�d�-�m}|V�;��	�`~׽�#��{#Y�Դo�������>F��U���)���&񗌔KMw��f�����fFҝ:���C} �CyLS�6C+�&�.�Ӽ�).�1􆄵����KC�ڊ����n����]X�2 ;�K%V���8��U��O����T��`{��U�f~�V�zd�(|����s[n�A���RH��b�������o��Y��#�-�JA�"+�TVF����5vy�b�r�,F~��GW!W�J��cs8�bp�sM��7M��
&L���-�~ߴ����!-��ɢ|ٜ��'a|]l/��n^Ш��
>`�.g{x����
e0g�����LR��4�	^��&;��@Y'yw���������K�?�����!��]����t ��^��H�:hJ=���o����=v��7/��<���ЅF'c9?brqje��(��0s�ied�&6�{Oɍh�����HԾ��Z7i������9�,��OO��P�I\2��Q�m��B/7I�U��/�f���t�)n�P�'D2���ߖF>`жjY��Ab��!ޒ�hlҐ��wU�7r�����Ϭ萕�[��ަ�9"Q����I�7�Lc���������)��R�f��M����2Y+H��Ss,Q��,���
@��υVB���4s�<*-b�U�6��&�)�qlާ(힏!u٠s"�����vxh��Μ)kG7�1A�����T��,<��I��K��W?��a� �X���O�u�ǃ`=���^锔�p^E�둝i�δ��;�
.�q2�P ��=��7k�4���_���L��%%�婝O��W�\�i�|��U���hIY��<-���ڊ�����ɱ
ۅ)L���8F�'%h�����8[���\d�Cu�$l�
���/��0Y���i����D'(���?��ھye[���H��In�a.����$E���K��(Q�hk�4�5~,B��653b�^����XO�!frTVvDNp=@s��5��Mcg�+�������A.mP�N��s��Ϯ`��Л�|H$`����VS3E���ńJ���ۅ^N+�|�2�T��
Ё�!�}JJ��'w�6~�. vFxnp6AĲ����9KokV��q��T�S�c)޽(C��ut�+�tA��ܻv�P��ϱ�$0�2��xM���pz�VĨ����T)x!�X���,��; ���䢽}��#c󓼨��i
��0����D�%7�����,3�
��S%D�Oq~{v�.��.u�J��^{���R�ڹ�.������sAYHy�k�-:c"��}K��gU.�ɜ��p�0\��wmR�+�B��l���2�>�Z�.bP�}��9؆-L���T��qjn�J�]D^� ���%qfnlhHU�
� ;zI��`m�IW�qO����fk�.��J��r�τ�W9�YL�N 	��8�\���.7B��W��Fq�B�|5_W�^cr���q��ٱ�Y_�c�Y�:W�vt� �z'1N���ஃ6 ��m�(�!��(�\������+�k4Ϣ����5T+-��!�cTr�Ā
*Y,V7�A6�S,r��iJ�-S}C}+���
L;m;�GU��MVV�l�,m����%��&�I80j\�Y�Vx�(��G�@8#�_��">��d��Z]��v����Z>*#Y��Q7����%��$�e��/�'��{9�wj;Is�n�=�7�����U,�(���(~t�T�� $Q)�>Y<"�s��^$@���>lXN�Fe�iX�_��-&09������Ҵ�ŸCN/Ç>�5 >�� �V��zu�dS[Rxİ�h�+|R{m�x.H�d��B������<�=:*����ZkjY7xP�T`��Xl������c�Y�nV~q	C0���)��^��t��*%͒e1|<�T���an�}D���cB�� �mu�jb~C����xx��P�sp� ��G�����RW�[��{��ʄ�F	��X�vP�Fs�-��ѤT�|f����C��d7��U�V-�}��I��\!k�>��Q�0ny�.��O/��<5��抣�QE�ؼP��n�c�68��;�N�R�us�G���_�r��|{� p�Ip�a&tg�+�3��Y���a󾺯�s٪xU+��o����P$���u-� ��v�0bF�:g���s�[��PCFta�E~��1^�hA�1���ګ�qG��K<r�`*�g[��?�f7b)���r)��3yke<�M{Фf(`nmA.i�#w����Q�o��,�#(�hN]�\�2;� ;2�j*�U�aoXX�����D`�B9&�u�{��x���Ģ��>N�~^�xE�m/�k��g�4�'��v&�	��@�����~1��_�J�z��YbJ(���A#۔e\8Ne+�T�[l�\E�]���Pt�2�f+�_�Q�Y$�/10_��=хھU�b�|en��h��k�Ӗ1Uq3��W���k(���+���2zT�Z^����Q�i�6ꔯ~��wֳ]��A�4n��A]�������/��:���կ�@�^�~�)S�V�����L/���|���뇋���j0���|��_�:�(�@�_`{�3�I�y(+�k*�ZP�>�>X��<�b�'���|+l�nz�ƶ�q� ,UdC1������	ߜ�w66�\�x�/9!�Y�)�׍��̛*ᛄ��9�>��v��9 70��%��#����	xr,�YP䙔_��U� �k�d]RU,C�γ?�=��$�hK������?y&�L!K� \fcU���x}b�!R�m~f:B���F���z�o�_��G�%�F@��Td�C\�[$s�`���עy���6n1A�'���}���^�蹅��)��=�Y�C�f�����P�i1S�w���,�$�F���� ��L%�����
&G�3��=��N���D��.�S���O6OR�yx�x��󘸒��$w���9^ƿ�q<�&�i��KR��.n]��yq#�m�O=�����]}h0�veW,H<{��\C�sr����7�יV}��b��HYy9,�0)���,'ehG�X���Yh���520`!�9u�@���]98��-������O?�6
�(CL5����M�֋Pa��J��}'l�;DwY����yߟ}�zNډ����ɖ�׳�[گ�5z|�9y��/1t���딚� `�_+y��)2�om1�RF$}���U�9��#lw��Y�DIc,��>������Ѣ��6H�[2b{;E��H��nA�'�{F�)o_fį�q�������$�T��!F=��N����ff���ώ��Џ�by .�A.��I5�cƃF��t���CX��]�'/�}c"�"{B���}�	i�������ɚ��؄�MXX[�����LH#ksu�oL���P�8ÁߧO1�6Ap�M�\9OP7��ce���v�/��nn��]�lO�=l������Ht�Y�u��Ɵ�\�<hмͭ )H����3�L����@����V7�Я��I~�����P�2z���l�������$X[����g�B$�ǟ��ZS�؏���L�X�7�n�y̫2U�L�>��\W�:�fSI`6?�i#�r��Sh�3KI��mH���ͤź��诧�f4�w:��ف�r����m�0������P����q�(O����y#Ȼ����y����?��8��:2؃�Jy�=ol�EV3#�SNThgA/3��?[\���T�TLKAp�B~��)�`�NtEd���Yߔ>��!�"��fWn�(����.���Ȋ�ѺԹ��GG�d���r-��~��k�㝔�C��u;�%1��K1���x��V"��^����G�'�v�828����iD��IB\��M/���޵G�.�,"��tn�X7�.�x�b�P��I�Ŏ�ed~�D�Vg�j��J�G��,�)8���kʲV7��4���m�},6��1��0%>R�!�����eꂕ��Z��#5�K������Ԧ
��j�n��'3��":��	�9����L� sZ��x2�]a�׃e��R�w�����[�i��=Vv����o�"����1u����7�L��KŒ1}�]��eO7gZ7�����]�W>C����-Ӯӭ��ھچ>�/��ˉ�)�mR�HFF!�Vb�~ա����g�9r,/F&���s���ĉ�m�W�W�D�ȡ���
s�R|7���U�����ӋȟT����'Cf�4~eM��=�ƞ��?����u�R��1ۜ��6��Qg-�5шC�Q�C���a��5����gc[s�O��`�R��Ӯ]	3ӬC8I�ф�\B��9��q�+ʜ17G z���QE�2D���_]yM��T�JXA�!�geXw긚�Ewj%��|��6eI����������̧���o�� B���|i�y��v��w��XӼJu�8��i|��8�k�bc�>���WC�O�qR�'sTg��l�Hc�Ձ;��q�ۯ]7�a�}'���S<����5�M����}s0����Jz3r���ԗ�\7���N��� ����l�R4���gfԔu��Jg�����IA V|�	�[W�;�$qĚTK+��Q�/Dy���nBZ{�����w��Z+Ԇ�z��exS��m�J5,�{�zYB��5��1��eå��H����\F�K����a�K��O�ニL�<�O���{���ܼ�W>�3��E�_)��en���zW�GT�����t$=��>}*���6�S{Z+?Kp#�bw����xͷVL|�
jM�3T[�,�[%���|�k`��URjyF���ɫ��������n��@����P榺	�9VV�ܴ���c��xFB��+#�=4G^�\�~g�-�gv�A�����Q�&������WS&��'�-��'�l4=�AK���uok��ǫkc�ܚ3(]�zN)�u�����R>��}V����s�����&�0b_Io�����U�,28��J���[��1e����Ϫ��?�a�U�8��UEn@b�W��~c90�`$R��%�5��Ss�v�1�`���z������6��)j��6@���05:U��ij��Px/��{C"��ԛ@V�ƄJ�r�J�~��[)�jA'�k�b��Y���i����Ȼ�Қ�yZ>�܊L��٘�5��J�Y3�zi]J��!eED���M����
��k��X
W�6�
a+:f���߼d]J� l���؇��[�z��ՙ�5�?��3���?���[�^��l�m_"}�a�9Ⲍ�h3f��Z޵V��]���.@O_�����o��E��Ka������P��*���Z-�6��`ˬ���m!הI1-���,Z��-x9��n:���`S{��Wa���=�wz�o�w�Z�	�D\�&�	9�%jǓxg����c��O����&s��K��m�`�#I�,�/��=J�M���%�
�!��n�mu�:%z���E�{SJ��]�m<k$���Lz�����ٔ!��9��\r��.5��%��d�HBL��^�r׋��a���<5<�D��n�pv��������%p�$� �G��~.�N��~.�@e�g�8W��k��ɚ\t��?�)I���d���6��Z��]��4Abϯ����C_^�xw���+z��Hg0_=c�̇���u��SC ��z�P�06n�I��� �\��鿸�,��)ÊZ~=��RCR@����+5*�[_M�8����$E:{�A���P)�R`�{�+4�� Π����+V�X=-�o�<k;Ģ4�^��Z�L#�
��2���1W*v;������-^�Gf_ono������Z��.��^�4,T-��T'���!����SKoS�L]��뒛�.!��������wJ���)�zT��B����/��{F���w�Z��Z{�dW�ͺ}#�A��0&a����b�2�Ѓ�q�gJ����q�	('>#�YX����Kq�8�~������g����V4g�w�t��=�Ԝs��g婵K�wѠ6?���>3p%���NC��W�9���j��Rɇ=z�
o9��P~����A���/=��kP'(f������p4��Z+�fP�N-�L苼��峒�0�8=��H�����ȦSR�56���7�g�3�9x�X���48a��e��$�%�{o��j!���%�6�I�G��_5�~� "\:�O�i��*/�̗�v�w�~b���	�!�򦌀�f��a�$
-*�&N�85��&�i��]��k�R��;��_P��s�g��3Q�ꦾ���Z*Ka��S�Pcq�;��g��wecv���⚅ˍ^�׸�q��6_IL��b���e�ҡ�?ե�Ⱦ�׉�LHw�ٌ������_���Mv���߭�3��y�>Uf�|S��s��J��������4{h$�T�r�_��Z��{�Mv�h�a{�	�'5Kj�Բ�-�6	)�����ׂ��}�2��`Q����k��(���7�aF�k���2�o��z��7>���I� ��gm^$5%O�7d5ߞ���XpF{��Tx F]ߔ���2���wޝ���.A���ŏ������A�Z����}�Ҩ������I�G9پύ*X�'����=Eʍ�2*s(+�1�F꒙[��T��	J�EIZ�%ww�{�b9�s�P"mJ.n>ߕ0�M�A�rU�mO�(�����/����n/��5$�l?���8�q�������'������ ip;��_u��#��2��lGX&�a�ww�9�m$��~s�x�w�k ��ƒ4ʯ	AY�kBd���P"�pULz�|ؓ��į�������Đ6s��#-~e���Vs��eB�t^�U�?W&9����|�9�n�L������k"�=�~әZ�P1f*b��t|-��fX;%����i�J��{7���[.(����@��,W�4�kb%��t�0[�#�CM�����^ݑy�V}VljYGR7������ҫ\��2�$�z��gLԴ�'nH�V*
I�ʅ]��-�U�9i����ы:�2��r6g,��H*��e��"�dф QZ�����oJ�ۓ��z�B�"�#��ӷ2�ʰ�t{BgeWbWf.�x�«��ɑ�:k����l�^�R��M/ƃ�bJ��\F	)?��� ,�M��E|�*��/'�Ԉxnnv0�mpgOVļ絗��-�����^��R9����:�lQ໔�}�`��*q�w|�qG��sj��fblt5U�@��Y�߈�%u`�"��CÔh�_�% +��u�#�#_}���N��~U�
�`g9��X����Wt��2��p�0����v��G����ڧ�X{3�Q���FK��F6�bx`��⢖�8>>ْ�W��4L�\hs��a���c�tw�{u½���^�,�c�ƭ��#�a���#�!m�==>UT"��MB���Ms8'[�p����}	ótC嶧�=o�|�yMi��ߎa:��oU}8�#fO��VLac�GQ��lե���-_l���J�S�X-.�"�^�Z��������N�Ў�R�9�Y%�q��*���H�=q�A��A��9�n��z��m�-�ۉ��k��(S��у"WA)P����:�@��������_W�2p��;�le�+�����C�6uv�O*[	�و���,�w5x�o��}(FY-T��Q����-H����rV�L�$���.�[�k���N��C��Ȥ�l�m�>��ΡP��p��à,7P_����V���������q� 2L,�� ,|½��@����\���aΐ�$��AČ�8|[ڕ�$h�?6hޗ�^,˜�v徤�BmKn�!��|�Y�>)������:�X��nj֗�{;jZ�wE��U���|g��9���S�i�����t���e�1Ce���D�֊���z��I��v�D�ɛR��䫊E�r������
od��Hc]��I�$�O�^���Lx�{�ea���y��B��C�oӚ�9���=t�������#Fw��t�\tK��� ���Q������P�h:χ�,����P�;��R�ڑ4�ݩ����4�	o�A&��r����e��o����F��X�� �T<ol�>��M ����EK�<�쓊QJ1%�1
��r�3�}��.s9�<#����D�Ø��� +W������$�%P��'��w�^���pCޘ� �w+ ����`�9�qг�Η=)�=���y\	n�`[D�}AÜwa�����a@����	�J�>��y5-��s�sfZ����2/u��.S<t�[��h����`�����d_��ծ��ڈ����BF�.%2�
eAdY`Đ��>�(}��3����b��R�5��;w7��k-��uL�mk��$?h��h5ebM�>��O�T|o�Ƙ��+S���\=���d��#�7\&*˼��;�2��޶��S�q���θ4Yґ>�]&�w��s�T��<��z�|hG��tX��u�<Ay���������Vl5��<G�l�F�:�C��^H�8��w�V�0��O�/A����pUϳ(P�0����痤��
��˰B�&D�W���W�w����Ӵ�I�ɳ�o4�W,�ۦ$K�ֹ,�F*�m�*�a
o�&߀�>�/��4��"m3��峰oТ����޼�4�8鉽P�Fa�T���U�,ь]��?u�m��M�L}��X!-�]_�ˬR�����G�%E��{t���ց�ۣɅ��n�``e��MSp�MM\B�x��'rsfX2q��E�,��8�
S�f�y8��Ɲ�q������sؔ�Q�eI<:'_��Cw*0��v�`�l�y8�p���UK��r���:G
|����')<�L��ei�Dy4�X�(��.��"�#���a39HK�	%KH�f���H&�{?�^
��U��1�#-ށ��]E���|sP�H�wd�q�����/����.��y�� 4������]$�B�h����gQj�z�������D�W�*%[�w���{'�t�G2L-I/x��*��I�R�J^�F������~'�݆Q����FN�EH�,�C�`y�D�����:?��2� ��r
`5z��8j�qL]��{�t����/� V`��y���[�>��{�V��)�,�v	׷�l�(�Z��Jm��4��˽��[�nke��9��tc�t9Of_�}8T�N]|6�<��Ĉ������g�$�2 
���9�\�ݮ3���\��-:21�OV���O_B92,H�#��]~��������'�T�k�a��5r��s	��dy��O�sª�U�h2Dؤ9?��
�I�M~/���
d����uOcܻ��7��>~�&K��$��sצTP+M�d�ӺCO@ +&�?CYڙ[9^u�Z
�_eܒ/X{;���^�y����AP@l��~=���̳�N^-��'�,j/g�  �����Q&�A��&0ŗ�0s��Ҍ��!�!UҺ�k!�]J(P4�� �W��$�k��D��^���q�@�G�W(�u֩��� X�y���Z�Tb���I��Fh!1m!|���v����LZe�z��� ͑RI��S?hm7���huml�@/�UaF�I�������3Y!�7kM��0 }Lw�3��3�
(Yr���Z��\�l��f!m���V� 3��^����L���kX��
Ӯ�Zt�V,|ߊ�P�,.jU��iU-���sò�΢u�����7�<<�ME����@�8��@� ]��f"���
�����ʰ�I~V�ՏL�Ab��ͭe��l̋����YXҊ�$�{�zpT|�|Bg��E�3���$L=�Q׼�I_ma�Ν�E��v-�+�L��/,G�-�8�rD(�1�t��>�9S���i����5�Mȋ��Z��S�\����>㗄\YC�Y;c���YI������'= �G}���o���k�<�2�D��x xl���v�}:�(��-_��X�bql���̄mTJ�LJx�}la#�Xh9�	y�]��$7^&	�s�2�դ��y\MVc�\X��lH��)v��`���j��(�..˩9�js�I�bA�5ҐS�����ʞ���z��D����0�oL���(~�z3H������@"��u:�z�� ���)��L&���Ǟ8I;��m� ��B@%'w��+ep�W�4���ׄʍ>~/̦t�����P����u�u��y.x��wh|e��m|ᱧ�#��bR%�Lmq_�_�.�MM	�v��-�h�m��{F3`lh[��G�з��TT�ǈg�b��F����)�[�C��{c<V}�~�APS��Z�e�9����E�Kӽe�Ո��<��11�*_g���B������D�7�ʏp ����sqM�&g�� wJ=�ܴP���uj=o���S�jGw�g�ϻ[�����g z:Ee�p)��M%�Os�6�#;�-���§=��>�Vc&�l�=?�ޮ�p���4�����Юák���R͎�s��[���n��m!t�d���(���(Щ{��At��恀q�A��� A_�c������?N�U3��ZIq[Gi������5rv9���m�H�"eũ�q��c���`F��K����.�h�п~Hy�ҫEbL�ܩGM��Č�Q7^�����_ (3/<�O�����<�A���UB��1���q��g�����C7mKPP�K�y^�AЪF߬�����j9��R,t<��?^'��נ���V��[%��0�1�5(r ^I������-��yd��E�ۭy�G@��4j�5
d��.Ä���<��iσ�n��Kc��YF�AO�$�Z�����Xs_t��MB)�l�oZ�{q��hu俼Uλ�4�f��W�͉��_e�J��V�l���y4bj6�����1�S;�. )_Ӝ�?�[-�c�()Q �������?����������juA�y��~������^b3�!*�@P�y�g5���_�zϴ��u�� }ﲿb�w�󠬣��*2k�c�[�f#���~�4x-6��A��{2p<�@�^��E�zG��Sv���!�:��Z�\�����C�a�l�.����Ѣ���Y�`#��uVl�L�}�?�V�����i�A^�hs�b@e(�6�`j�Re)ܶ{riݣ���	:�b�h�՟@^�rs>��}v�T��]]�▬}���h-ڣ�����b �  j�%ѩ�ԡ�� J?a���IT<d��ۓZg>�gW�}��4.���/�:8���i�2�������������sc�^2������g��v�vt�����
u�mǌJ�۴<%z�p��vP�|U�/�t�p�HLm��~�Y�f9�;���k\;#T`�R�s��彘Բ&����Z��Hd`�KZ�`<����~s �hbg�4����86K�$,��&pK⣟ �-��_%D�Ѳ�*t�hj֫\���I�}#��p��pN�ը���^u�V0ף��S��u�7峒,��7r���3�-�֦v#�v�?\	�^�v<I��~*B���)�/K_��L���s=�sB�;��k���y��".���_��l�`�F$J/r��M��2�����TU�u��o۴�ɲ�ImV���ފ.'�(K��a]��d�|����:��X:��,��T��T�"��[�kd�ȍ���O������|�xm��o���`�i��'���O�4�^c���C�~�2띨�����?9�U��z,�s�Z#�9�
n�-h*�������q��,�@�8���Ԟ� �$n�A�(N�����/�r|"8ySp	U&�?�:&8;@]@CW1�ml��
"�xhxCLv����W6�n^&�䱣�*�]�����r������+��"��8���${��Sǌ����4��R�E�� z��[G�p��J��5���Ǹ�������IM���u�ƍ�_��4�i�{�v���]5����{��ߎo�.d���J`��X�]�;T�n���Ӱ�Lg����`D1Xh��Fׇ������CV���X[#��a�c0�}�kz���0o�sP(n�G��,��;�v��l�kDې��gʌ�Z���/2��Xn��ב�;��F�k}
_� �j��{`��Lo���x-�|r�_�VvL�[l�2�5qˠ^�F�z>4T\Y:�+�1P�0�t�Ռ�}�s�����W���qG�_�s�o|��ԥdv�V�z��Ӧ6�L�����q�+Z/�6L�Tڟ~�l��Q��!��\>�f�,���fi������>�S�p!VF���Ct�+���&�pj�,��+N���4�?��X��*Vg�>���3�->�t��	��m����Ҳ[q�G��S7�
Z�f�VQ���N-�+A��Ls$��k���[��Я���T�~u�Mo�:�i��!��Ib�ӧ]�=HC~VF]"[�� 0B�z��KM��M^�]I��ey����FuֈvU߬W��i.��)��8�_<����itpgoYD0����|Àv�;����Fb�d��a&(��1l�Z�tSJ�䷛���B��O����1��}{܊bX:m�T�q��^*
��Z�<$T�� �=3*�;�UwO��f�U.G:gy��z=\��c��qB�p��|�]�0mwڅW���T$J����&A���WY~���	���V�/G�}�7(Q�^_Uap����)��TtKݼ��	߭A3���Y���IH!��+��}9�
=��;үH�y��b��/ɨ2��\{�gQ$/��]�-�����<����������&MG8��L�GO���e�[��Q2Q�L�
p[���*1L�0�(��?5nS�ןH�@�ڎ�L�6�3�҉�{l�wk��`P�_T����]�g�B^
�>�\�W)�4���wz��X�g1��'�#O�n�� m5���n�������t����^T-gӵ˞�'���=�9m;�����%w:e����3� լ��3����f������Oq�S��ơ�Zf��I��k7���%�������F���T����u���3���6���;�@�e�)I��Ž�����X!cImpz�#���_��}���ş�+}n"!L���Y��a"�F(G ���-A���~����1,�O%��%P0/���� �A�[��n��SS�2{U�H�;*��l�!:,1	)�c�y'U��>w3�7�+e#L?n6�S3���ۧ��)���z+m+�	�b��)ݢ��1+\�v�.��b%�j��3�׿H�L��G��F�&u�Jiz}�A�dR[sYYK&�0�?����O��:���^�ב�p^yk���`���t�n��h
� �8�_Y ^	_?|�<�h(�w>��/{�}RЁXܴ}��#���2�q�J���*�M�P:�D�g�����E�m���za �n��uo!v��b�MA=N����c%Nm�TM<q 6O��؃�8Z"`��������Xw_X�R�[�S��Y�s>%~�(_�"�u�����)f�D�Ѯ:`��oPFϟ�q�AJzu�~��StXK<%C���kl-V�̇5�i���Y���V=�F��׿7*���tc-����j;\�0+rQ�Vo����m�������Be��K��fΑ5z��(�u�?��Ԕ��e���UD������+�_1��Ge���Q�D���ΰ���|��u��&�5ح��Q�T�2��bԚ��n!��/&^�o[�pU�_/�5`n9|�\E���⩵�?u�*�̃���0~�L�t�;�k�u�L�YJ�q�+B|�݈��	lw�����k97Sc�G��S�B/5�ba��p
z6���-ʦ���}I�X����GD
��~�F=�����9ь����*a5�ʄ�;J^Mז		k�C�p󌿯����ZMG�m��{��U ���feq9+���Ƹ��|��Sq�mI�V��Ζ�N^��Iܛ�!�(u��԰z)�ǫ����5�n-0�A��*Ә��k4ƻ>
tʆ���6>���\)�1`��	�%.}�+��̽(��ϸV&Iݩ�g�����&�KJ�ڻ��4/ �5��	-�`����&�/�'�γ�W�p42�?��.1�оp/ֶ{ٸzP(��qBn}1&K[ן��滞Y�Z��*�&���!f�/�H���h���#�$X�&@�����=b�7��P����/q.&�0�AKGH�GT۟Kd2�r�d*��,��Tf�fk��:�Kq�Pzظ���]�M�05�`���f]I���Γ,�X����AS���8�L�%�{���uw�>7%�2`gy[��k���ᱺ1^|��B�=�@J�-Q�~�ѣ�>S�ƴ�����V���p�,a��o�.��#$��l����N�բF%�*XNnk�n���Z/�[�S�)	���GS*��"��_�N�N�X�U]������1�YjBON7KBL����
,�Pwm�V�(B\���WL�o*�����~v�ʡ�(s*�C29Za�'@� u}���Je�h�W�<AQ��VZC��= !����vy<�֜9k��m]��iO��d��:څK ����}��/КP�X��6MГ�f+��՗ä��Bʳ^�+���)k�0;�׼�p�i�.����S:���h?�j��	Wܽ��j�R�������	Z�yiv�`t�PΕ):PrC��f�jw��t����G������R�BR������r�s8�=�NN*<�j�{sA���~�	Dtl^�DB�z �j��#�\<ܨ��,/jj#�$.;�h��G$M~�EL�(7yBul������aݤ��!�f�R��
��˷�3	��T/�����1���|ׯ@�}��Q.crx�����Nǃq�!!��lh��p��$iEDq�T����\�~���_�q�v���W"R~����_!S
1��D�(�Sn�{H�ӟ�܆���)蚲x��*0�kg�B���j�%���5�`>;#(�� ��E�[GE��}ã�(�GPA��.��T�K�CTPRIi�f�n�k���f(��70�9��}�k�,\�g��������{�"�����	HI;8A��yfa=Щ�Y$ku�6ZN���f:�T�,��^=9׍�ekїM�qBٿj}&�LV��ք�oi�4��{�>t�^i3qo�������E�Z�ߖ�v�ݠe�~�A&~�K�Ӂ"�@�_���g�r.�êY��a������h!%<������J�@��2���ӷ���B��d���T�܁F�8�he/
F@�ad��e�����Ѳ���Y�RtC��B@R8w4RZ&��)�`�l���޲�=���?�[�a���9&����j���K�����5�
�._�K��/����G9:Nbǩd�W��㬯p� �����JC*�v�0�9Csq����-��~@�Q`�C`�"�ʲ��%�K��,�6�=�v*�V"��"�i%�{�"�ŁP
�fA}�S��QhlL��}pLv��xӴ�zݎÅV��,�oQ��k��~;\o�
����o��
�P��K�����l��
�Q:�<n5�&�B���������<|ĕ�4�C?n ˅�i�
���������l_L�"G}5�4�ԠJs�����Ƿ_�3����a��	Q8��J_*��Mp��er|OR�z2���OS�+�6��Y B����:���ҽ*���cX³��*K�qՓ +���>}��]�PI���]c|<����%i ��sCI�r양�rG˘F()+�L�U�f��a�����T�ڊ��k�� ��O(�A��[���e/��o3����s�X�*�^�~��Z���u�d��x����^�����9*K�+��l�k�������wO�5��OV��eZ��D(���8>���?����kۣ~�%c �g2zw{��U0�-��2띴�کP%�h)�.�2[����ݠ��rn��c{��n�5�2�mɤԧN�d�,�z����W !2`�w,�Z�z�],���s���]�T�hu�p{�h��LpI#�y��`�::�B2�5��<w�	��'dg��y���f�>&�:M��+��M�g�Jz����y�+U�X|��|�f7�{cY&�Co0嫥��2Ն���7m��r�L������@���+���`����*2=Y�R�s/��[�\����]y���2�$����%r�\�8�C��{]4�����_��.����Tl��E�?�t��kRT����M9��QT�٠��ց�9l`d}S���3�&)uF~;��f�s棓�8�~�j]ʝ�,r)L������ƞ6���5���ƮR�˫sG��W��P,]m� ��$W̿#B��"���H|�4�l|B��'��>��f7�G�+�S��d�z�+l+v�V��Zb`�i3Υ_����]���_��ת0[���:]��3�~�X�1K�7Ɩ�j���'�e�(��/3�Y��q��J�-Ixٝ�,*�Ƨ�`�$���c+��#�Z'@k�,!�az[,}`KT�E�nXQ����x�-&Ma�Y%���̓Zs�4v���,��̍(rV�5N%gؓY�5M��!ߜڛs��{�q�-ľ|���D%Ax�O�<׿�������w]5qK���q4�eTdW��gʆv�hޱ�����&��$y+m=B�yػ��h�qiFR}Z��xA����5�_� ��9��Y��g}{N���̢��ʊ��i��X�i��pt5rl�In�?x(/@u���:|����!�}�W�[y�Lbg�/Wxk%�w�����̚�,a����-S��.0��tR�]�;��S�\�D�"J�ܩ�Mv��؍�����I$.
���rdؖ�q��$�{�25�b��KG,���r��q+��3��<�fX��^1�L��|�O.�
�mq���J�6�2ލO�SA>E-,��F�-�~|�q����.)P)[ٳz����D!@f����m]���  ��i'`D:z���k�D}��a���prF�h��<����/��|��'�I�+N�DSؽ���Ʒ+�Li���!����۽)<���^'�
%��ɝ�yǎ3��O�P������P�'�Jn�Š���&YvjQ�c+}���T�sp	��:�������6����-yr���8/B����-�0PG){ �C�5fɛl!���+��vګ�j&"��|�����#��K���#Z�y���i�L�W��� ��t�5\�y�i�K����n �j7���� �ѧ�ӧ���ܘ���d�'�x�f��$�P�{S�"�X�#5A"h>@���z�����T��(���R�vv�L)�lٽ�d�$�.k�3.!���(��.`�c���X:{l)%������ӎz2���޲T4�#U#i#"��?:*=,��aj ���G*6��:��51G<S�
Ƴ�7�WI�^vJO���+ը\���9	8JwĿ)���p{������,p�	c��v��j*�,ٷs�M�=�y�5�M=�.��.n�6��ql��-�Oo4Y� \Ĺu�,7[~<z?J�&�� ��
Nh�AJ��\v�̦Z<�;�8���]Ł��@�[ۻ�
����ӓ�i�\���1�ffi䡻��`�(7�,�OD��l��썹� �v&k���L��g�h>�3z�����U�#K���;�B�W	�5�&��Q�1��S54��,�3<Ogx>��!�6�m�?�=�L$��鶔5>{�Ǝv��(/f;�b�Ł�+�xA�q�/Td}*�ZH|�<X�	?�a>�z��N�c��~q��%O����&C�0^Q�N8�	
td!������PH5N&���q&��ᏪFU	�&�XS�jZj�H�ko����.}&I*���!MjQح	y�:��&�a`�l�,�1��G���d���4S1,,TJ��	�*E!����&�J�"�E�NF����P�S��%	5��7�v�Ŋ"ڢg����6�ǡ�y��˒_Y�t-����6ˣ˨�(>�pE��G�7Cw�-�����[b�*ܧG���3����;>%�MA�(z�I��/�E��P��|qP�}=�I�9��ҥx�!�X�[U�On��ѭz�gK{j�P��U��Ðwg}�qɝ>:�Ď�8{}Nx��N
��� F8�8�ꚨ��(=�Q��u�$� ���+���~YG�����#���ߵ�w8`�4��5SҒ���c��׾���u�"MJ�0����!�.�nȇ� �Y�^1�/�G��y��^��8���w#��ӹ��T�;��ϙ���dE﯌���ȅs
XTНB�u�l���/dq�zi����فI@��͛O-)�Px�W�P�4��[�K-��i�?7��_�TUBp\��N ����$��(>)]��m�0]%�,;���SE�R�Y$�G����T8u�'��f��(�fĐ��mGL�5�01��}Z��f/jxw^zȼ�$@�|x!:>�č!�f�O�z*�L���3�q��N�!sy �*z�	{�Y#͡:�u����<�,k�+�>kmԭ��7��2/�#������.�s#ObA�6��o@�.,�E{��1[ �f�YXO��ɖ֨��Aw��Ŭ�#<p���W�R�s����A�9�قKL,��NE .!�l��w@x抭����Ԟ�(>r��s �爙�� ��8q����\9j#�{6͚���2�z XZ�斛���_�L��M x(���xo��@������W6�Tp�6K�Iܢ۟��Z�BJi0Ӆ�ղ��"tֺ:��<�ϓ81�?������"3�ݚ��uKCeMI��*����N������>YZ�2V�?����N�%� <����VO��)��N	�7��S���p3�����q�L<s���G��r����^���`Y����|��i��yX|��C���(P���O�|�\�Ê:6��ѭ$v���e��6H(�d2~�u�Bz[,��QU� �B
��*$�a���n?̷=�0�%; �f��74�E��d8@�Lm��}�N?��k.xRT�HsX:��1/^�XR.�mz�.C����;"G?�E�Nx�C��Y@b-�%�p��oŐ����a3T�J��� `�!^(�\����½��Ul�����mȱB��q6�n���P��X:�	���B�U;�/F� ;f�*�c��}޺��𱒜�5d���8���8����&;)�CY/���q ���
~oki#��8�X_����M��F5z�j��3y��g���{��]QU5���kM��d�Z���m��?B; �@���={�8|�"G3B	&�\�_�q9	�ڧ룸'�X�^J_�����U>��7+8E9�Zk�/��>b6H�m�]��=G�M���O�z��JӔ/��=��7��`�}13�ؖ�*<���0h._֜�"D4��H�O�병<�-+ ��[�s��Q�N ,L~j�2[�"��58�M4G�׈���Bl��>%���ӭc�^�_J'rd��ۭ����6jQ��H6���G��,J����`���fg��F<��ī��Z�R���&�+�\���&�9�
j����<,I��s�o��N������ڭ�(|����޽
�������~���Q�Y<_��պPb��h ���ص Gzh�Tqf�\�)��\��a!�n����G:�h��守iD��������Z(��(��*z/����:�?u"5�:���$'ݓM�p��k��UN�w��>e�H̀��r2,���0���P�vl�]C�}��vyB�iz����`/or&�7[�y:hwS�y�Ez!*�\N�dU�ܗ�o^&��,��~5G�ァ�ݽ���Bi��i�Ç���M�ʞ��|�Օ�����JS���}R,�Te,v*^�R�D�a��^V/������֥I����+s!:*ʳ�-\�3@I�6Ә��ЍzvwO��>]z"�y���{��z��h��:w�na�S橣��x��Jck��D�S�x���d�����+}U�Sq(��3����R�6�q)liE/����p�VZcܺU�OaǑX?�Z���k� j�2�08U&0���j�O �p�*��}p��̣Q����Fk���W-2O@�H<3}����Zޖ��{��O�),V^���wy�j���Îp f8MPVv%K(�E�2�tI�`��c��I�����p�Hdn�#�ي����4k@kN��z28'����Ie£��� ���Zah��I ������=�}�i�.�� δZq��T�E�i���iO�L�t.�h�H��eqz)C�l�.��t`n:L��X*�TE֙aH�8��M�*ѡmi��ӕŅ̷��jd��@����\��D�%S�4�ſ�z�����CR�����$�O�.<}�q�Q���8�K��<��}[��QC���d��\�80Z=�F]��G/#;�׾�ح�8�30.0������v�'��3�2n�t��V����+�p��.'P�Acf��DPrr�+2�D��'��z�!����S��.vKRBpyHn���:U���-D�A���wu�h�i�n]V�|���z���A1���WZs�������o6��ѐg�"|���.��jY����B�A�y�~��N���ϱ�CEs��~"�@y��?��L%��\��T��*��w,�f�D��)J
����� �<��
S.�M��85�:-�ХD�7�9��R��W�� �w����L��p��I�}�
+Vחɫ�g�b��נ!2ܒ~uw�bv[�bG���qN����s~i�W��jD���G���_��ò@�b�~F��}����r�ۧ=�#:�%"׍�g��L'�����c��b�u��x�7�_�
�47�PIZ~�]�`�*��R�co��P�*b�wO4����a���#�)Mv���;�k{�fzU�k˜�ᬭ���!�|�S��������f�v��c���h(C��������j���Җ�����퇿n� �C�-Ȼ�_�k�hsŷ�b��#�U)��-Aq0� ɽA�#J}�1r���=���@�u��)2F|����h}'�/{��)�_������Hb�a� ���X���� �]���d��r���I.S��1`>��r���*��^�Px�ƚT����| )3;�/��O�N��+����*홑C%L�h�|�z���ik��<�W����r�Z^�=氁|H���R��a���?���~G��C$�_ߥ�Q����\�9s�%ǅ�Z3�~S0eUG��۹//`�[�������E�ݯ��|��S�#|v���iKS '$Ee�A��h�K�#�-��!.�C��¯�t���E�,?���=�W4��>��R
����RI�b����R�epB���K��)�����Z�w ���
S�-��l��N�,�
ue�難��20~���a�e�`���$�^"L���T���������a @��

�ឩ�w�hd���M������!/���s�?^S��P08��\[��r���Z�}߼M��|
����q���RdnY"�[q@��q��T�������B�Ru9��x���J��y��v ��/v���ԖP�\�B��� �t���Tyj�b~Lw~ORm��2�z<ų��e$��� � iW��c��I�V6��A���Y�R�4��%,�A�Χ��6�Zs�~���K,y�}�]+�a��Y�& �̷Z?4�W����$h�x���N��!wG�c�Ɓ�H{C}eT%�}��R���n�I�[,α�9�<��K0�@Si@\||WC�i�s��d���j��Sa��E,	�ʼ��v�'���Y��}yq�>�M!d+y#P@7��s��T���%���X<V3"��z����4�A�P<��q-����o�6)����>�|��|�ф<������їp���b�	��-a4�SX)�}-晢�(t���m��Ed�P4�	9f���eK(|RL����bĔ���F�]W�ࢧ;�}#�-a���	ҊoŘOwNލsh�?4j:V̟Pb��`��P�y�+c�b���H[��'��}�\���NKi�4)��F~�$����z�̟'Š��c���l�{�����:=�p���N;q���,5��0��p�OL� �L�y��������!%v3����kSV�g�I{��ʰ	���u-N�3���j,��O�M�,����9�$�X2q��+���h���9�Z���l�ՠ�{W�Cb�\?Lw���nd��!_����ً�ڻ�d�.���G���X��Cf���aӝ���k����S=W�y2<��7�J����vcG=z�������Ԛ�Q1���%`����c+}{~7�6=��Ge��+��_��o�(�r�rS̰!�y�6�����b�,c�p���|��«�ˀ;xh�щ���Y�6Ou�E�-�ͽ��(�� �����:X�4��%���i_�|r$���7�Q����D�T��6jnK�*S�Z��;݊��= �y�֯�X�+w�ͻ �#��={p/cz5�oXiN��@����_��d�D~=*�=�%����ɩ	.9$HK��}��/֤�l\�5`lǪ��Q�9jڏ�f+CrP~3�o�]bsQ��y\�gQ�ف6�5��I#Ji��cY�VC�ʱ�Z��Z�lFӜ� \kuc�\�����wT�n]�׼�z�W2�T=���ϵ=e�؈�F�-�`�S�[�L�.w8g4:���<����O���ܴ�0,�Q��D'�fB)�e0_��*EEEB����9�YSmg��c@���xQ������y��*�D�����P��&$_����L���L!�J\<�B,/����]1W�Co����2���nT��C!'ޜE��b��-��b�U)�%�.ӌ���)1�h�FR�~M�y��(�b9-S^�v��O�A��_v�T	������{�2�l#5�����B���˓=�^�丌���Z@��S_˥�eg�o���_}�-p����|$�>����<I�K�7���k�he��&_��{�!А�Y�xa�iU��2 wC��;b>�r�s����Le��-��ݓ�y�(�_�e�� e�L-�TnH�����z�ד���
aE�,��k��n""�FA
̓p-���?1�_��(�9�r1w��i� W�Q�`Z�Į]s� ��E���\� *)�B5 ���C�h.�$����l�\�4O������E�EI�Eb���8͹'=�'HE����"Z&3�&�ёbS !@n/�@���t�
J,~���f- ����u�� �z��f@ڗ�nsqg�c�2��� s�������+��TtM]CE��������a�λkFS;j\R�+�HIW���>�%Y�b!�m������z�M,�c�^��N3��B(h���ʹQ�Y���~s/S�&�S�=Uh[�I;z� we�g�ف{>�ҲO(.��T�*u{����ϙ�yj�Y��2`�B�>�&�R�ck׶��sX�TliA E�P���S}Z(
8��4砄����<-�c_�|<Y��%����G��T]��؅uǡgpd��ݧU�E�wjc��'�ι����#a�<��X�'�$XN�&�4�8�[� �X���n#������rEm�_[I���3�t"KU@�6R��]������n�HI�8�0`�|�q6~.��[�8�O���VF�c�ae�RT2�jh�7���\�0��uf̀���e�u7�ϗ��A�t���ւ�+�pR$�ʥĐ^��A��9��t���\�{�2�h�G�Luv��2�/^ty=߲l�'!X:������׊���H�U%oW.�n�=Г<X��nUQ(��*^tٴ��J�༼��Fe��W�08ja�y��O�K.-�;����s�N�� ��Ԯm�?Z��}�2���A���<u_�su�0XxH/@P�nZn��ӥ<t��{>Hr|W�@�0��nH�nxOo���>����(�����TwiƗl\��O2���֕m�B���gX�:w��l��D�|��D�zd�I�4�V���&���H��O�$�yZ^<Bo(���g�����\��@ة�=����p�J��O�T��2ܪ��V����N���E�RY �/�ٿ ;;�fou�^�z���bkK��N25;;�	�X3�U���#�5�+`ܱ5��+�W���F
�7��Q�Zۘ���7ߕ�Yb��N>Nt;�\�r�u��HL�zU\��,�<f�@0��=Y�δ�r�I��|,���)��L �8�9� ��⤰�����1�Fw�"��I���5ϔ�P�-��K6�T�u��X79���&��U��U3�O�VcPn�ٟ�۟�@��w�VQ�;���sz�XX�R�-�F�5;ީ��t�_��C���nF��/��|ѕ�=ةe�^�w�D������?O Ǳ�/W���%��!�ð��~ �o8����:[c.=�}KG����h<̈���t^Fq�c�����"w�c�[KY��/����������s�'�iD=����Sy�Q^9�n2M��сJ���������m����>S�.QZsY	����,G��֊�|�;b�=]-���T�b[�0��0�RX�ʰ�A��ی��޾w����\%ɲ�')���7�
��@�&-/����6O���Kv H�xR��o�\S�1ބJk��}��B^�L��Y�Th�騰�'�'�dMi���Wʐ(u��&�$���JS�fJ�ҝG�����SYLe� �T[��s0t��C4a��vw_�m��!˂��W �`Gi%7�2dQl����ԉ$����@���Cko�z�șy�s����W�b��~��;n��3��� �ߥ����L��ô���X�!�I%�3�8{�1]M��.�|C��O�@~e�B��I0����ed`��Ȟ)�b���88����QӼ��~�QN��n5�ޝ�ThA�(RV�,��^�qP���W���R'?58LS V��"��@���Hgb�O'M��RȠ��+�yY����:k�Ļ�~js����Ȧ�su�;�v�ف�l�3<�}�yi���*�:�*b�i�d���p:�ȷ�'��$���U;�|����T64LC@�g�8{5�=_��h�E/�JB�u�������=����G>V�j"}Z�.xG`oD�-m+
t$#���������S�>��>y1����dLR��|>���<�#T���h�H �	�����~�ӧ蕈�2��%�j��/3Ŝ����0�yŪ٪�c��4'1۷�n�61*�,��i��c8�A"�v��p�����2���EW�
���G��bB��C�;�����	: ��Ju�����x���G��FA"��i�z��wN��zNN�g�fo��
���-|U����6�g��Xr�⃮qCc����~r]��i��<p���<� Ή��:��S��nټ�o�6 ArE�� ��I�M�?Dh>�T\f�S���)9!Y\D#ra��dy����|o�#�R�:�Rj�3q�E�	ъ(�gY�BIW��!!\y�	�PV�6���6���MZ���Y�R�J7$eb�Kx�4�q)b0tK�bc�d6]9�{n�g�ơRG���W�t��/���IL4����I�3�lf����W@��ϴ9�GWkx<�I�����:k`��0��О�{�2���m�W������P��� 5��>Ԙ�;��SMa�u���O���0��޴�}xݶ�� ˺u����[��L��q����$�|���71bc�Ů��x��x�#���n��O�8֛`�?y����^Z�����L�$u������q������7|_����\�Ƣ��(�I����+�~��R�6#k.�s���qC����>�F�ܬ�g�F�G{�;?�,�v"�	9hdÖ+@O@l�U!�R�\�>�7���c��J�}[Ǜ��{����;�Иj�P���[̲��I�.�!  hLԒM�r�)�Ch�O��PȋN\H�i���l�T�qF�8��+~����L+c�����/+|z�
D@�U�P"�`�=~X�4�(�)���r5�}� j�:��*=��U����QI�>���G�~��
��b�Ο�)`o�ħ�[�μ_����p�LC�36��N�h��58�(�x�ڕ5�peq�ݪ5v}�4 0��^=0)�F])5���絿��db��������+��u��Qx��Vf)~W��4#U0F��te�p�J:�6��f�K�Tf�H�;�\�����b-�b�6�K�#� ��nF,���٪�p�m{[�e ��q��s-�M�^#�Q����g��ϧj�n�U?>5��Rl��	�4FO�ᵵʪ��M���KŢ�L��^�2]�T'ya��9�,`}'��8���E�3w<���T���W�V8��rXG� ��/Іve�Sz*��5�N�x���q��(�N�*{��Ry��M�%	�{�E����P�78�����G.C�r�g��(�{�	TH��
`���]����{̕U���5D
��DRr"�+Dz����w"��?��5�G��Gk�Q���u}���^��}UX�����q���R;�iI��9�xhB�D�&4��'G�EG�*�'��N��L��'�+���;BdR�D**Gu8���EHN��]���?��}|3��x��Q���I$f8�V�	���	�}���x9��a�����q�Mh�E���"�f�钔*��Y����
݅=ۢ_S���):wL�֪���ejD�~�d{��~t��������l�)p���li��Z՛����-�T�3�_�	d'`��R�˞J3����I)|�-�c�I����������/R�q�s�����B����N�Y*�N��_O�b�������?�I�~�1RY��� ����m`��g,4g��}�0t�謙}R���n��]sYb��n�,���CD�H�r0_������ɛO��]��B��u3���k�s��s���3����Ƚ����P	����Z$�T�Nі���T-����C�L�#Ϭh�G:L2�$�b@=CJ�}�v���V��˜��Ψ��,G��?��pv	h�����߷s)l8�z̢��P��y|��~74�-�k�e|G;[���W�x��z��KGC?fQ�"r2�
�R�n�-�R�m���f �����= T�|=R��%黅Gԉ�b�֊H,�1���ق4�������sJ�",7�uDh���j;áZ<�B�@�3�W�#M�h{P�E+� �V�l�N$1���,ӰNq�m��A��x0��;WY5��{��ʨ"����Ș�L�DP���U�s���J�(+�PV�=�C�b���˯<yX-��-ĘuKz��te.�((�&>���{)��K{1Io{#�0,S޲h��� d�o'�� ���$�ƀm`�����!�'F��;I� +Ņ��~nS�bZ�5��(�ڟ�.j�Q����?g�	V�ϫ�[p����"�3��_����"���v�J0�]��Q�w�t���9	�W%v��#�(�/Ei&�q��)�i����0Dȧ������aO�3�8���۲M���[�r�;�������L��<�|�4ϧ�Y�}I�jօ���Z���Ή�� ɽ��+��UI=mͻ�o�^���������l�r�g������\�ԅ�ۜ�L�S�0Y�SIl;� ��O=�p�T�vǞT���rph��OAf^B��4l�Ot�t�?L�M�Wa�2�"�Z+`�a��}���4����v:8�cA3�����V_��gfg��2�:���"�m��qꙎ/U�� �6g�I�ڏ��锇ʿ���$�j�T�vntt�v�3��:D�5��-�XI��\I���C��E��N��B2���%�]!�J1�rN�슥mb�%�~I���0�Y?Q4mm�Z�]�^�fbz�d��F�ٷN*��.�N����]i�h:74\џ��}���g�6�Pa����;��1;/��LR30���x
�?�T�E k� h),z4L��Zǵ���=/?^k�I��>�;٢Ƞ(�f`h��
�A�u�2K̆�K�DEEÞP��P�3\'h]�� ?l��>�μK4��[�z<�o���V��X=�|q��z�h���������g��xR��q����n�_-���E��q}��4�2#�Z�#��eK{=�h��=@|Ɇ�Q�S|�P��|�\T�u�����i-�vp(�n�	�gRcȭzfw�{؟+�-^�E��kʹ�||���8ǉsv�e���|��{��9Q�f�� ��I}���%��Uʃ|�s-���l1�p���w_�d䶱��8���F`�K�AO�u�ΰ�?y#��ܜ�`���,ex��h���hkn�� 距�JdK~�2��t_����|Y�
l��|��v��!!���������?�3<l�?�!a6D4��&x'DF0���Y$�wp0=-�9S2C�������ɫWihlD��̭M�����x�.W�԰�<,Gon҇4�����cn>�JN�#�ȶ��O^�I��W����
"V�'r�'�"�,y?@e?	)����XU�D%YŸ�Qp�ؓܐ6�H��qJ�_��l��[1t�:�ͼ�+;�lt�v�v\! ��M����!�F	cǽ��2t���`���8�����Y��r#�/w�Ō���q��Ź,Gڇ���j��	�F�/��V����;�/�ˀ�|�Ds {O���-@��h㮖��k�xR��R3�r~��W�.I�4���{��i�'�=�iX�`Z���=��LUT�Hc.�:{A�.������ׄ�l���^�U�r����W�7�M��2�J��z/|YZ��F��h4h��
�\�2�GU��V�j�"RRRi,,,2<�Č���	lw���;� L�v�>鈑�H
����?�z4��h��֘�d ��b���L������&�m�3f>-)?�*��٠�W��ܜ����ν�Y`5G�K�z�xC2�-J�nE�OM�a��5adj�е�w��7�Ae����)���|�X-^/2�}�П}�QV�G�(B���q�b��6޿�f��{moC�����]���R�ߧ�!�V��R��_yfcl>��,S��}��g�x�D"-��8����l.����x�귆�B�\���.�<�}����/�&�T���t
pg����LLL����#�H�q[H���.z���gT�:�ҥ�1
��]kW �"~WRb��}�9_��3S�����.�Wy^�劖�����Y��y��ҥ���n$�U����J�6ЈQQQD�;+**��{�Z$�������
��#�����!g�)�ħo��%���$麂�Z:�hO�÷:^V��H"�Vu� Ӕ��5[�R�����@]��`5"`�!ӻ�X���n�8�4����?[����8��L5���V��n����������%f����t�#�AL(^7�C!pk�sQ��c�z������S'�"��^�FD��塎���W?�.��c�q�p��{�o�׮Sy���i�@x�*ig.��GOV�7�E^�Nƕ~�&�Q��)�p�q��������T��&777�"4|�J�'65X���j?ʻH{���Y�e�xWkM�n�����_�p� $����!�`0��,���}gº.0��kO�V	��̱�-tV��$�[/*�J4F��Y�ս-J0&��M�i�p\���+��Jy���! +�:����P�T:r9-�^�l0���ɖG������;���׶��*$W��H��qwX�E�1Ͽ��J��1��X�j��K�{�(-�ݹ��?���C��ф���gJ��� �UN��_���lsqh^
yJ#tC=5D.}��3BZiʽ9���������3�r��"��^Z"�F 
��.fH9�*A�-���މ�x,��g��Vjv <D��4�������*=�'��;蜼63u���EIFn�����W_����`oK椧AM��}���h�x��C��g��V-ti��.P�8[����B �'TUU�������X��>`ͧp��C��!��F[�$����?�R)Ӧ��6U*:��:�ӧ[9e�<Y������.�]����%�t�k���`bN����]B���O��E��/�Y�Z���L�S�\�~����r�lÐa|,8�Q���?��z�N�=�3F����Uɚ�yMS�&0��
0�(
��_�~��1��*:c��4�62&�4	eM�B�)��7��S�iqd
i�R�������:�yԹS�d}��sr���m�bP�'6zed�1]�I4_��vRTS#��q��%w`��|$/�_BQ�7����gHV�8��f`��Y�!���I �t�{*�'���iB���"�'M���g:K}q�l̷�ׁT : �G��e;˕��Y������!�вWR3^�_��|���=k�/-�z ��ے�����2g[|�{<���kk;�����&����&�z߼/X5�;ԩƆ�=����n���615�i-�/]�Ѝ�.M��jc�#��}w5��:�������'�T�_�&��v]4�:��L�;�`�̤�O��Zo�nL�� #��|�>95!�FN�Lԡ����6n�Wv2�u���1���C���y0���m�,�V&�P�����z����n\*L*.�\��>388�W���e��{{���T[� E�q�m!�R���ZqQ�a��,����j�~��e����7�s�7�w�@w&[|��r5$~��q Y�}�E���e���QaF�ncUNV٥4\A�Ɩ��u�0�-""bUO�����Jz�w�Η�6\���Б�N]���շ�u߿��erV�" �#%B�Lgw��0��r��W=����{%R\����^��O)$0.d�7�:��l�-RNA!�����I�ko{zz���4���f����#��(�J��� Tt�GƄ5F��}�	��Gcyi�?��Vio��Z���
��9Y�����4��yGi@�7&,�K=4�};=��ߵWm"M'����Qh9�D���c<���u�����1Wܑ�m2(<~��Qz���M5�$%$��i������oՂ�̵�K�i 	J�=j�����A�8�*4l$�����@�e�x�0~�1߉z��#"Ybb+׵�xP�����	�ZX��Ht�J*y�@$��z�t^
�mZ��xA  �!����J*Z)#c� �iX��^-��s��`�]D��������z�]�44��ñ��Cn��I�9��Վ���^ /����a�o��`�l�z��6)H�/?���f����z'-�o$�ɭ���R#��
1�rphz�����L����g��7�f~�% ��u����X��������I(�[��.�f\��wƶ�}}}n�;ȝ#�<-����Qy��РZl��J�ų=:�z�E��Lrb�Y�������Ttt(!��;g^x�ޟ����HyFV<C�K�b���%!Lw�D���s�Ѵ�r^P� �T�޽�!`�ehx�c�/���an��i��GNS�O���Ó=,o�dO	귄:�7!t�.��&D�֣j$���y���J��Ptp�l�yyw[Z[	#q���6��[���w��!X],��Ȏ/R<�,r�j:L�S2�V��m���<�������N�!�~��WPP �;444����Y�s�F�^���~������t��KJ��!jg���;GHS��V(��o\]���P��5���Wg��KKgdg�����̯C�	�%���*WF(�6���ޟU̒TS���q]t��Z�+,�/tFq2�H~|߂��q����5��񇌁��R8Q�cz�S����v5
���)��xy���:����1�0|͢�&�������fm1��a�!	ߥ�
@y�V;����^�ם��@���
��溍$��C8�4�K|]�BM\���o` |����Ռ�Q��EC?�yϛ�-;�F� SRR�@0EA����L�����2��p�Êi%?��n�!���!��}5%Bx��b�����ɷT�O��d��������z��F+8�І�Q�aaaY��؇��X�|�_1�c``�.��d�r��^��.P8�%��������Ei���|A
bLղOKs5�� �8Z�\�F�� �
��?d�Ks�7�,tl4���]�I��7�ފn�_� "`��w�̓�xGlO�Xh9�-D���6��uK�Է�k;쬤�4Z�l��k$' N��lqq�h�6��Ҭ����	M�!��65�����(�L[����㝩����֏D�xPa����:�\N;�05���GI�f��V�tyF��\�95�#�8���@�K��>�s��+�;�����)�I��d�rs�cKV����Z����a^.��m�r%�B+�a�j�sii�[�����W �6���.2���=���l��RaIq"��;�G�O��x~�58�d+"�%�U��? hM�M���볝A&������y���+r��o�O��f-˺��P���UD��Fo��k�=����p,3s��Wܨ���˳���W�lI��
��0-�U�p~�8i�Lg||�P}���恣��1pq���Z}s�$��[Z[g�wS���%��;+��s�w�-�;bڥ��R�N7�,}�Y�X�:v���8�����ӹs�׏�+�����,���箋h�1Z���Q��'im�y�t�uZ��C��qCI'��=<&������-��*i��4�gҰf�L#�����@B�����ўX$����R��ܷc�߾47�3{�I��u5{r��AߟS��ZiIC����TEho7����q����_��kw�i)��N�f�������k��W}��HQ��R��⥉tiB(�	=� �NP�R���AzQ ��[$�WCI��?'��_�b)�0sΞ]�g�=3.=�Qt�!dwx-����P��{r5��"��j�|�AX����Yj�������kV���k�e�),X_`�Z4Ғ��ѐ��t���ĝ�`�^�����ƾ	V�����_��2��j��>:
��Ž;1�6���V=�\�ճ�G+� �5a�e��Y]]]k�������c���1�7 E��0��*@�gK�e�"h���_�
G�4�4�
�����Wbz+����P���:ry�9�������7u_n�f�	�H�L"���v-������1(((�S3Lz�� ~�<�c��oXj�������r����yS�|�=f�*�����k���/�l��7�9�W��^(Wc�&�U��#�+�����`o7!��46�̵��w}�����pU���L������xP���*-���!��,�%���`U�C[�v�~�p�"��<��^s��3%���[PO8�^�{٩����/��<�ޟ^�k�Ř�z��S�f_�����]oy{\lz8�/:�:-]zQ�|}:55!T���ƖY�Gy�A�=�C��+�ڔ�i�Q��	�lO̮����M�m��>�lK�_�P�Y��+�J��5�܂���3N���GX�h�)o����<C#҅�X����b�go��˗!AɖC��ۛ5��嗩g��uI�}�x�����YO��a�L�7�4*�4�LA⿂�7�����,�`f_�PW�ќ�b�����2�OF�>��- Z_KI�d�>9�a�j���H}y��!$���+O�0���N��A�۲��0�p42A,WVnoM�+-��зρ¨-�q��9�d�����M9`��-�����
O��o/Pt�F^���m圣ߴLX�52�,��e�k���Z��:z.F�iatA�4�z �Sz*��?��r�]�)���@�Ԟ�~���ߣ�m��%�����ޮ����f�/; �#��e�������2�a���o�^{x,��΅<P�n��a{��~���&�\P7�������H������)8�*�LsJ�鱺S�~YsH���K�k�!1uw�i��n�ѵS��_𳷺NgU-9����AMAM e��U]ӥO�Ԓ���P[���V�����M��N3?ۉ���>}��*+ua���+y�ֶ���h����kc��nY�Fvn�f�-�Llf��+�7�����^� ��v�����_:�p���bO�!|"oG���t���{�M�C'�qg�-�p�m��kB.�}�u�����</�R�,s��0�o��T%�� /Z1���L��VJ�!�`u1W���U���`Y�b��]`�_.�a[��o����5# Ă��	�G�bw��.C�6��8L��MFM�y��&&� �TH-�h�ͽ*&��!��ÙL͢������Y�n��:�u}�ׄ��RZ�4�, "�u,T�55��ĆR������_Ň[�h����9Q�C�\�wP�w�c������:<����|�t������B�����[��� �N�_������c����K��=STYfi׭�X��jv:�z�r)M:���tz�!��lU�A�÷����.[�v���e��k���84�0lU�0��穝ƴ���?d�A��
�tH`�(�_����튒4�I��k�� :rb�ѷ�ǽY�H�L� ��e&����|d!��.
�p���J�ysWˮ��PY��Px���P/���Kq_n��~3@n��~N��pM6�#+g{�[ʝ�%kS�+^�t'�4F*�?4��1ʠ)�w�c����!:��� �yI�0LA� �x�K�Q\�.����Т��b%��������p�6y�`v_�R�ߦs����V�5;D�,'t��]! ��FV��D5���p�0�/4����fQ���+�@��M�A�
�[�x�iS��2ɾл�RQ��(zѱ}LD���D�Cs����� ϩ�mhg1����T���hy�׋�L`��_n�k�Y�0����S�k��e�����:K��?��4珔$�F5;0�/���2��PG2�L�ݓJ�����*?����dz����cA��ThX�R7�VD\\���锝��R�ؿ��N��7�Z4C��p��W���j����Y>`��;�{GEE�i�-��݋� ����6ճt��~�~��l�ĩ�[o���`57dr)X�5��2���� �!��J�܍����]�C�$�����iW�����q�^���zp��co�e�(������*q�R1g'M��+v�ۊ��3|����yNj�^���U�������M��\ܖ��i���޻��+!�?�b�ʰ�����
�e�T��0������P7U�PԀXT�����N�q�{�a��EipL������)��m�̎�����	��0��'��PN�}�e�nxBk���29���Ė������o�SH�++������N��E��aEĦW�Z-�sS_N4\,)��}��=J&��U�:f�RGE����q &��.�q��bZZ>�5�v���Y�!Q��V�t����M耢õ�� ;9�����E4�
�blY�~a����5Y��<VO��[�c۴!_���,��!�Mf]�-	<���7lM�T�O�67 �RU��)CrT�7{�1R�#r��B *�����d�:��Ӓx�rv��A��x�n�����ܱ)�	'�V�$��*p�2B﵋;w[(�
�� h�g�d��篘��#���
~�X�Qp:����i�%N\n������]yꂥ�+���f��<!g	?��_\�*�_��8�~4Q��4#9���Ju橇-����>h�PI�Z�Xi��M/��"Z�]�0a��Z)WU�n^�?��|�k?�"����Ȍ8=������_��C�F"	��ڪ����~pLx�zu^Ҁ�ia��o��s�Y�,e�u��5_��FDc����h�2d�����b����U����'$$��]��De�wi�A'��a	���,W�UGZ
]�� l�@q��[���H�6�j�]sEkUS��Y��*2,��a.W%�����}W�0=}��:*����P�EN����y]���r���an��K&��DG����zZ��uſ� 7V���+��k�q��a��&��l&��,rw�\�e�?��?e�-KDe�r	0v/�ey����ݩp&��+T��K
��	��>��<
��� Z/�����:t`^�!�c'v���+��a��Z�����a"���g�T�
A+���5�U��� 3�;���ȗ�]yz�+D`Հ�|��{�l�1J 7�����U-�hgH;60�\s=�ͫ�o�Ǝ7X�39�},M+��P������E������ڛ�6����K�a��J��+����]��a#�/�ve�@�X�R�%�v�����K�L���^�I�����f"f�?��Z�1�M��sHc�>X��w~7� �������Y^�,]�:���0$�ɋk�K���<셦U��U���r������k�ʉU�O�ʕ��y�tT���F��O��}s�ln���駖�}����Y�n����\a���L��7��\��(��������xC"�ߜ����	��2ߚ.f����S_֍�s\<����\|�� ��s��(	l���8u=�No��wb����T����D�Vk�[P�sMm���9��v&�� r�}��N���H��%_Q^��x�H��$�r�|� |�j���4 7���'��P�ng�e�<0�m��;�$л _+J��t�=z{G�r%�W}�h�5=�~�v�:�Q0�t���چ�2>��|	y��'�ז� �xd<1��^Gf��㺟zT��ps΋���4�]�[�F�$/�t��Yk�Yn2zp�������ad��/�n�~���S�NKƬ�zz#7��d���
�O��1��b��,ru�H�	�����Lb@��-�8fZwK��Z����7����䥝�F/�cW�%i�ZP9�O���'��dV<2�v`ș�e�a�@hC�qX�U*+�Ž�� T�U�����=����fM[m�G����r�:w,{r�yM8�N&>5E �$�ڡ�Tף������0��mVQ��:�@J�af��碑��<]��c��S�I�zCe�W�^��^bl��E�*-n��66���0�w>�iS�����n�O�2�l�ܬ�����jQ�f��3�T�i�A�cD|�,��AWx#���t#��r`�I�b�w[`4�;��J��������KG�(&6Z���f�c８i�K�#Lؕ
~$ ��i�wa��ûK? ˑ.h��5r�T�# �h�nF�s�2\EUG]_�ү��������^a::�U֛G�v��;�#b-�ӑl�n1q.�ހ�]°1�۝=�Ym|�J���B��!���A�$ک�~������ݾ6��K{4Ӥv���4\nE��9��1���-}JV�!�H���0�b>=v3u"�[�DU9��G����߭�k:�^�G���e�
�U~��0�b~Zn�?}-����:.�32�,i�	�F����������+�-��� 3�m�e�R�>+A~�'IL�X 4OL��!Y������/%��]���3+b����TS����&S4G�]ec��E�$�6Ǭ`�<��6l�+����Y�ܺ���u�D=>��3��G@�����\�� ntc���9����K!D+lp{�M.�Bd�ڕT��]��CƼ��e�x�������4�n��PZ��*�JZ(�T�X��U��LF���[Qn��noo����a��Ҍ�әO\~7������\:w���~$�9-�)n���b.2A�U��i�6����~\x�dJX|��h�����O��r�xC�p�m�`4�g����;W0�G�֮2����}}��㉭�� ݅#7�  ����$�;YR�y��ҫ���Q5��oH�C����R�z�J� ��"A��5�o
�9�� �kk�@'ehఠMh��������=�@�����eU�~}�۪�h��z�y�X��G��U5뷭O@����~�����,�c��s��k��/����
��/�c�i(��
pPWR����zMO�:] iOw,�ۣ!�ܱ�.K���k�A�ځg9�J4ɋ�*�?C�	��c�g��:��6��(XE&���8l~@�!gF� c.S�o�_>|BU3w�w��k�9�(ɡ��*X\�)5�� 6��ѩ�#JJJ05����>}�"��.���0KW;��-�Gm,� S�-{�Hi��~��ӑ� �h��*J��|��,+��+�B��z��q�?�g7n\·0L�?5����-��=�p�}v�m%��7����~u:Z��J,��)�w���eAN�-�x���[�+DFGGZ���埍�һ8����n�{�}����t��S����|�=@�i����K�v�4������-�k�h�.���%�ɽ�}G]��J3��4 �-�g��5!f����v/�i�@> 7�E����e�vs��!6�?���s?x�,�W�}(D]�d|��@���nȭ�ʹ��\I�($LR�z�3��
�q��D欿��23�J�`���ڡ?%<��H�d��6�i� �r�*a��o�*.U@j�� R S�(���%�FC��a��Csꦰ�G���4fOXp��xl�~�K���3�K\��<� �Y�ʖ,�:�ƶ%����u%?�z�Ԏ�]'�@�P�!}]3)��ߩH�s�kcAY���<��	L$f:qqu
��F��3��_K��-$;�3�"w�����~oP����^� y6��ϲ|>)5�}����nʚ@�(���+��pF�D-#�]Ẋa��,r"�"Y,��I�0G�����%���ՃmHy�n)�i�G�l;@6�-�(��(�n����X���#n<O<&%U�=�RX0��ǄΠ��2 gU��&畠h�u{ �˖����2���Jl�Y��̘L=tK�	���C���w�6�&w������U!�z�_�??x?v�Q�>*L±�6�X�	�yuE�;%1����G��&6h.m�����#���P��uF��lm���h-�=Wr��dZ�l��(��HN�)��9	-WçW�P+��Z�n'+�8�)�:u�Ss-�S�G�J\�w�7�K��nў��s%�Œ�����Ɍ��~�7n21�^_��3�N|��炃��e�Lԝ��hz'd1?�gØ����G��'�>;�([�&6���]_ǔl���$���םb)#���$�~iYvy'�����0mĲ^��K�(u��������Hi���)�T ӇP�X3�X�^��'w5��G�y��r��e|��qg�0j�(w9Y�+�0���c���z�U9�{�E!V!Й�Y,�`w��j����O:4��1\e�� ���9�&[��4�vxt��)#X��;N���0a��
�� ��]s	)|����c�
�#ŀ����9j7���R\\tH�@���"Wҹf�|w�0 ��l���+��v]v��V�Q.al�W�<]g��G�ɇ��7�� hRqw(�$��� ���$'7䩲n��s360��H�?�u���k�30�aW�x$�~C-�8bwʽ�(�a�ފ�1���7�h@V�,�0Z���PpGs��,��Z)22(B]fg|ް2�`���V���ќ��C��t��h���Xb��d�p�� A~���_]�줫��b���`�@g���4l7�of���rD�h;�#���������Hӏ��zu�aY���P���~0;]d����&�~�):��{tA�8��^��oa}Nwd6��,{�s̮
�Ж96>k`{D����S�w�'W�|2�+���Pa]t0�)��ˢh�+3�[@�-���J�@�-(�i\܇�R��5��[P5{b�vLb�dx�����3������6/��֧Y~Ű���o��<�ϸ�s���?�6�����d;�Z�V>l��;��2 �h�Q_�mbF�@y�;�o/	�n/��"��|w���1��N�+� �GN`���9�?�G��uc�N�2��S��W(���`َ���`�q���{٥Y$�I��< ����۳,�6�|q��Z9.�B�y���/ѻ�}��r����,���ᝉ�<� ���aN�oO�E�=N=- 5�)'�ey���<K�(��r⇛=LX�{����^�l���j�V�Wy��Z ���N��^|¼t��Z�tD#ٽ���������En��f!%�O]��$c��H�@�D��I�_t�f��ᆽ�$\Bá��ʀ�It]s��ܼ�z����A�s���	,�sP[z�H�Q�m�g��}u���$�@9a�OxZBv�މ�p�����bBa��J%iE�(i���F�8al���a
1����%�zxw,�7ғ�N�!�F��5u����O,����h�^5��r,'��1�\>/��+S�3�mS揞��"B�#��2�-��י*�,};/��M�h&,ՕW
T�W�f��+,i��X|��Ny�PAy����\Ш�MY���|���X~khl����o.4H�mF'���=�u��Z1���πK�V!LeiX؈yE��!F���p�8�mX���[�W%��Gq:��m�)R�m%tB��>��W�ͻ�,����n�z��%��U�e��SɌ�а�쇥M�h�x�v"ʶ���ڤp��Ao�9??lb���,�|&;�#ް�J|�i=�}�i��	�7?G?Բ)9����X�3WU���1��q5g�d��� &���?t�G��?�֫W
vG�r�DM���<)���|3�, �%�46d*�_-
�p��J��2=�b�} #�� ��2�YGC���y�/N�0Gh^�@��<�4+�<�7�]O����Ϗ��mJ=�WWXCM��1W����fF/$T�"�����S��7x��bZ0��m��%jjN������+K�r��X��Ht�&�,d ��9����g���q<1ȇ�X��pȋ�����J���_>�(Y1���?>C�:M�7����jqiIM��y�������ӧM`�Y*Mt� ��a[ꡚ���]���u��G�>�"���ϐ�RRRX����t�40��5���15eX��KSSS|=�N��i"������n�;3S��8y`ķ���أ�� ���5�4��n5ӹ���_�����ٳg��l�:2������S6=����Z�za��vz|DD|*�:����S�:����K.�@�� ���[�>�������J��ƍPu�:������:������?I�.ZR�`�UG��.�R���~�q/�g�Mx�`N�L ����y�u@ ��@RV?���l�׬��g�bb�	f�v��E�K\э������3VL�:��~����b�VC������!�İ�Ț�z`�4�����z�,��4�!|~�:�����K�����6�x9c�����bN���~:FM�+��kk�D`����[�/2K����M����©{䔎ԅ'�G�q��jWhd��Em��`]C֧i���f�����!XX%�*T]P��ǿ�t�����w��8�^.�Y0r��/|�;<b�o1ٍ��j{����B����sB���j�g�ɮ��n��p
/���t��yPHy��=�ɯ�Ŝ�:}����o�pW�g���l����X��eo �&�����K&I-�ŕ۞[8Z3Ʈ�P��)ϧd$E�!�2!d�0|����M�����1�1?N�h�:u�c��!Ë4�={��'��}j����w�+����ZX<S�k����Hj4�����9�_��O��������8���{<]�H��p1gVhu���M�gB��F��=�-��M	�N���>�4b8�������/�.���7�f��_�`aN�U��i�Z�c5z=�t��!�u�bX�g)�\/�b]���l�\/�#��
�u�2��.?�=@d��u�<�J�����~(o	�]����!jM+�B\wLmR���#���Ko�_b���vcR2��^��P��?����-����]�8�(��%��F�b��'�&�a��ȔY_��Q�QT����qXѷ2���#[j��+�m�U�aK��Iݤ�@XG+�2D�?����"�ǔ6y�P�;>�>�e�q�ћs�#������z��Ϊ
�˘�-��+K����76�0�������5p���Oh)�~����S�AE9""RN|4Y�#����!�Va�LPm#ɍ&���ݱ��!�,�r�x��Ҫ�6�������~v��};6��d`R"�}b�\6��*�a\��O�������\;�����9u=�؃[n;�k�n��_�;849��V�����7�/��]o��γ h��G�cG�c��R�����5�2VK
T���;xMh�ph/q�����xF�,�ak������d�#FЫ5�����Ԟ͘c���qbw�DzZ5�v��k<�������.���\��9&�&@���ϾS�,j��g(�/��q��L`0/QO�&񣍻��S�(Et0(+����ȣ�q&z����~�`;h��̖*+�F����|�掤F�: }��i�x�Ğf��gi�Z9Br�u^S�{~K^�d���":״�-�ՖM�=/z��=����Sox�f�;ƙ��KD�|�&�
���s%f�f�a��h�҉�&_���nrm��?Oh����kg��8E��a���JgS����$���7�5��|�n�ۃF����tN��ċ����Y�p�~�\����1m̔(3��L6*�����_m�E(q�y�6�OT��lc5}\ kM�Sw�J�o��I4�o�#E�� w���w�E֎��w��d� �Eҏ�9�s�c��$F[�G�'�z��ŠE�g��3��9����X��ar\W(�I9���)�/��329���<�5E(FoL��'����Rp����b�nSw��a���Ԛ*q��w���/(,Q  �'��ߵ.�jK�(#.gj���:Sv��N�!{]q0J��w�����u��c���q{�`�e���N��byJ�\(;u��c(W����qE����9:��ތib�J��\�|՟9$tt����|驒��ѥK���ۨ`]�8�S�8�;[�;�g�є��:�(�,����B��T�nl���ұ�}�ٮ�{��J=f������/#��/C�����~c����(G�׽QCw�/�Q�in�Xɨ��h�i��!3��1�G����H��SR�#ם��z��&���&Oc3-?��)����q\�͗�h,��N׀2�4���B�L�����/�Ϫj��C�0���/cK��������\Y*�x��K��HG?>��zzh����ūV�P�b�y���[V��bg�4T	���: "���a��.�J�Z�a9$Rz���.#��<��>=�s�Z�n�i(��/,t��G�����w��r6���OX���f�ע;r$�9B۳x��`3YqԸ�Ui �)���?(;�/���62�.�G�������	Fꚛ��4�L�L�H���yN^�+V���og�d�k =$�h��z���M]U���T,(�&��O�?s!�<�>g��tȚ"2�o��'.�U�aaCL~��[߻�����0�6�q%jʔc}��≧���L
���G �QҜf)��ŷ�Jo�lԌ��i���.:DS�8�җ��\8,,���@'�:܉i��.��$��ѧ�����!*F�Ŗy�j��k�̈��TV�޳���c��+���ruԲ�s�<@1K��J&��>omz��R/����O^]gp[�>�<���e�����ܡ�8^j�ZN�y�xn��c���Ԡg��H�����X��~�qK�I��:U�w,�$,��'m͹����n~�'���\��7��Ὼ x��ɾmk%�S�y?�J�wN�[�z�MZo�;B����K��zA��狠�r���H�ִL����:c�B�7��Ew���*��S�^�wiI-}��HE������[.��x�_�?��j� x�_vM���Ϗ2�c���W�ڛ� p��Rc��������:!yU��Ax���K�Q�����yhP�jj������K`a*�{���
�t)ʺ�����\&��/��u�gqG9�S~� ��1	#�>�;�^����#.�L�F޷�L6�Չ����i`����.��@��6?�!�X1��P��5�{%t#3+3�N�gd��)����墜"�R
CB�W���3l����P�Ӳ��xmyQ~J�-�BǮO�<��s�y9���MK���k��������l���f~��ɇ|/�����˾��\k�1���'�w9�Ȥi)�u�h��%����r[:�G�c��aRt%�6��w��$�ܓ���q4E��5D.��*�8h[޼�� 4 h����ђLʋ������.�+�����[$��&og�PN)ޗ9lq��3��f�a���m���j�k���.!R<�`��g�M��ɼ��L*ng�-_LCX�שc�npL���{/���rc�km���zU����.����M��Dr��IO���:c�,�z8��}�c%[��m}ֵ䏶?��{p����+e<􃳂m�e���V�S'�-�PZ�3�%p���N��y��ژD�"s�ƹ ah���%�z3�~���X��t<J��gU�a������g��O)�ѫ��]�W��QuM8�l�����6���+n���zp3[��25�D�u�V���� <�i.q�m����Tf
h�d�z&�q�������Z�	��M�7��n��ϋF>��'8��[�����~�x�Xau ��/<34���J\nߊ��;����J�7w��ᴿ�à�u�GP���^�2�u�Q9Yّ����7 ���R�gMUy6���lL��Iq� ���Of~d#Sq,��=B��z��aw޼�'4����ڡ09�#�e�2w��u.d�v:�F��Ε.����Vy��0�Á۸{㍯��3d��5�%1��gv*ѳd�B�OA�mN��ǡy�:�Nɽ�%��.�Ƃ��O�˼P����Չ'�_[b&Q�6g�w���m2|yt��d;Y�1���ҁ+��ʠ ��g_��y�}��Qx�p�������9���qV[fɢP����(ܞSRw�W"�9�eE�Po���9'9����V��k`Z�����h��x����A˱}�����D���a�|��I\�����Q���6�>�>]]1|�uN
�k	����ѿ����  *t�!�L�ֽA)��Z�X���uPl�ס����!WV_HI`C���_�$N���������U���݉�4��Gh	ҷj	߇KЀ�p[eX��ߎc�׍�K�Nm�%,��TjBN���� Uee'x_��#?���'�X�Nf����n��>���+6�S�ί� �Ѓ�SlxJ ����-�����?��X��u��B�Dq�R����ӚQ�,��[$���,�,տ'�m (l�v�A�Ӣg���kJm�\�D��d��3�C��f�[�?���a���Z��W��H+�j��7�����f�����$�+�+���s��8��z�)���������9�';l�Q ^���%��4Yi�PY՛�� ǹ,x�;�<].*��1�𳔝��Ű���T�=��F�����̹��W~��u1L��L��J{�8�%9��p	Զ� �T�Ib�,��i�K���.�,���}f#� ��j�f5���ؘ������	�4�Yei2�=���N�_��[V�(Z���b諙Ug7��J��lE2dh�[̈Ғ:uF���	Alt#ot���9�Pq���M�3c��b�G&4~W~�3?D��P7�1?����M���ǯ����9Z�t�J�S�9ӌ�]��' ����� NFZ�!�Â_K�P��:MϨ�2����0Q�XRX�,*,Ļ�ϫv�CK2a�����.����Ȩ:���	��[�~Z�~���Ӵ)uНB��ܼw'W;V�l���N���2�S������T�{y]Y(]���2�r��7{�}�(�3�TK&������ �$ZZFfl�2�O�0[>ۯ�w����FZ��ӋL���4:�����Wz ���U���hr��B�ׅ��N�'+k���0;5�¨��!�e�_�0�&�c�@Э]�_-4�F)~��@��bJū�U��|�L1|��%o��rA��ae�H��k}��gs�9��K�E����{k+��oNC���L�tD �%����8]�:�?���mr��V=hes���%H�N�ܜP�x�`�J-�O :��44}C�7��
Z�f�Ų�H3��fծֽ���HyI[/�ٲ��t޸���>0O{|�6AKYd(���K�@5��j�ң%{�O���](�6.LC�,��z`��R�U�Bsfa[�Q��EeMk�iO���!�$����7����|�A�z��z��ͫ�\��-\�����:Lf�8l�����H.�}ć4480�B�e5�f�ori�z�TA7��ɾ/�f�Z"���j���U�5q�C�P̡o#�u	(e'��ߣM|��m/ޯ$���S�ݠNܞ��Po�r�����TDc���ω\���V2��i����[K��v60�|�M���e<��g�6��գ3n�	]9ȋ�B�譧B���4>Ḋڀ�;Hç>��V�Z<�p{2�xptxГ�`k㫢J��~O��Zd�X�l���GpH�~��6T��
F=_HP�q�ؘ=;#|�Ժ�� X��
�KͶ���H�"��d/S̅L6��¯���Um˚��BS�n9�`���Y��RtPl����yM(�x_"����� ��ǤQ޾���RJ�	�8�zLo������'��&�Ͽ�Okj�p1.���������!���$m�P��kQk�!p�rhY�/���做�Y�E�lV364�3�%�$RM��]9��>���Wl�ayh[L�D|���b@����/#�z^F��.5�D�E�@�^LwC<����~	Ջo�STu����O_�Z�y\��ҭ ����r�d�TPAiOtQa�d,�u����ox8��҅J<;�7���	��BmG7rB�>q�3x'�#?��VW��uS�}S�7�q}�"^�o�����h�j*K͋�7��N>����`��jB:r*�Iގ�t�Xޒ�ox=���W�dT��/E4Y��JK�g����cCIiE�V0V��'`��z٣t� �;Y=��E�{���%326�j��w�&����:A��s�c��B�v.�`/�~.������>3ut��(آ^-�����"{5���O�k�߈ S�SGcq�P�����Õ��-�m{⃱� O,r��}f0/0��a� ۈ�^edn��+/JA���)�q��c=�8v�N��DXSS�DE	�������_)v��z�mo�����4��('�iQ��kz��� ��C���s�LE���r���br0�JuC��\{@���~;S�<����#kkkP��I+Q��vg�&�,���8�U���^Z9ʀ��]<"%��sGz�y�)�p���L�37�㔇j�#��j�"� `f�s��~Nr�}�(�����9υ��ܞA��ɩ� ;�e�P
m��,LQ.�����L���e�k�`=��\��cL�`�>��/O�G�_�:,4�߲��U�A�w�{�J�Nqhct8|϶��e�����긕�W������$.�fI����T77ٌ�=[^���&2d���w7� �,�	T�C@5�w1�:��G73�p����6�<i�w��׵%�6{Sw�T��8RN��Y�Zd��w�i��$������_x�z��t�LZ��B�8�cSSM����4�TJ����R�΂Y�/�� ˮt�5������lU VJI� 3�?�Ҹ`�z�L�v�U1�X�Y.[*���:���Ϊ]=$;z��A(�Qd���>j��V�M\+B�!�q��3��'�����ka̺�<��.�`K��Xg��q���������in��kd6ʹ����"����v���o_��Ӭ�"6e�3w�+綒��$W�0e�bN�;tNh�n
j\�1����oؐ��PR��h���e:5��Ú+�БԞ������ϸ�����A����
4�� ��D~5�>����!`�w�ʕPVڷ�,���L�\��m�m�RK���ճ��fz}][f�\@�JqI!�.(~�$A���)�� �fS��SQ�f-�Ƽ B��bk74���}m���Fn���7۩�4�u�@�V��Ե׬��6�~�*���_�犏Ss�?�,_e
4i�Y��+�2��@-3%~�-l$T},��l8�r��I�^�=BU�:C�u��Smm.�w�瑱�/e��7yҿ�I\�t_�/LZ��p W�,�l�Q{�)�EP�N���x�%�c�����oF�n�[�%/��y+�'�,��p���(3N�l�_?:!{4vښ���i����kB�7�� ��̰�*#�n����@ܺ�0����o�O��bߊ���WĈ-�]�5M�#�6�Z��ݦ��#��'-�Պ�Vz�󣏫��L�\@��Jn�ϡ�Tt�F�wW���W�6 �_y} �[����B�x��� /�wpN}��f�(O@��5��s[ӯ�B��&���}xX�$���T�4#c����Ẽ'(���&0�,F�����1�@l��Q�Ԇ��`9)�Q�Y���57߯珤�Ov�>��Vj��K^��Zl��oV�&�)\�`���"l��ky�ܜ�$C�Ceޙ�^O�Ϯ �.\�).�t�=n' �F��	���s#
P�\s���M�#,6�� �O)·��ty�[���-%E��Iӗ=�����Z��g>��Â�^��8���r=ӆ�>B���,D�����3e�����.��8�V2��d�#s�S�1���u��ΰ�C͋����;�aCc�T� �!��
�M�=$��S��������R�ƋC��W�f���ke]��}��S��yn��5㉌��?%�&�(+���R^"z E������6��3�2�7�
�"����I���|ҕ��8��7�Ys�:s����:1�/���7-<gvO�v�� YD,�t�����W젉�/" �����a[e 5R�]�� ?��
��D���
k-�WG哃)�!_?ݣM.`~�=�e�<L+�Z�9��({�Uy�T/sOÌ�N�T��4���eA�(��x�FX����I�<��qr���/��y�`�j����xpa�A��۫�qX�"JK9:Q�+bذ���.3� ��4�E=��V���v��F�z�K�>��#�0�R�bt|���,!Ҭ+��7�1���.	�S�������C�]��g������FN�-_�1RpU��1��o�k��zg�y6ۇ�ֵ+�c��[���Y��0��rD�xT�Z~�67��A�D(�'�>?�t^}��l�����<����E&�XJ����I{�/#�֣jDr�,ذ׫>\���p:����H�J��-���7�� ����3IM��(����`�̬�J���r���{,��z��xp�����ΞQ9�)�WW�yi��Ƈgp����0��\�G�gb�ڵ�;���W��cۈx5c�~�v�}�lP�������qR�y�w��u������R'�:!�g���QVy�/�~ݬ8|��L]
~ɡ"�,��]����S�K�[�t��\��=�nm��3�F*�i�
\�{��j�A~�F�4D}�����:`�y���1�JA���=��7n��#2|�>��sk�?��N���DX��A>|u����;�F牡e�	wY2_ `���A1Yӟ3�G�/���'N	
�����k��x�MCꔕ��> �>}?q3
��~���h���zy]�d�~������G"�Jg�`b0������--,��;뤾�e8�C~*N<���addds�e�h�_F�g���z��?1�Dm:�  _ 8��ܡ��{��J�R�G&��a��*�=�i�!�^�M�%���3�8�,T���Ւ"�s�<�}qcC[ꬕfc
��J�&��R�G�Ŀn �:CX0�y���l��c߯�K��X�X.�&��"O#2��G�%?��Ӗ�����57O��~�|T���F��7�G�Ё��%�~{^܀����ڨ<���-0kXJ�O5�M��u\m�۬���|%��b���:9d/P��X�p�� k�2� 8?X�M��3��L����&�ik��R�����Wןؓ��<N�3�B7�ϯ��x���<d�Թ \uY
t*��<�"�-�-a/StY��n|Xn�G�d�����+�{}}�7A�y5�x�Y]�|�,m	��>Z���/x�%�䤻O�s	�ܳ��ǍٱXR��V�y���U�����P�A鼦���5�����Q,oN��W����_�<���<�������@���i����g���Wn]��_:OU{�o����ЫH����
�*�.\�iiQR��n��6 � �ݡHw�t�t�Hwljҹ�t����Ͻ��9�Q���ff�����Y3�1<,?�L���b��Y����8_		���y����|�i��V	c�n=������2�$��ݹ���{�;�0�J���u�� G��[�������o�!@ۯX�gm�H%�(>�_=�!�?M ��-a�k��⇴��Q��������,�p��N��������f>ϓ�4E"Z�4Xy��¯�ޞ(������N�{���W�O��7��3��<z��G�ׁ�M%������\�$���[@*��惺�L~&h��V���~��dɀ���ٙ���������z�iN�e |c�q~<���6]gg���ݹ��0k��d�W�v���ᰝu?P���,/��:dI�~��_�`���6��i�����ʊ�u��E����"�ճ1"�y��G%M�'����ɘ�2oY���7�ܞ�9
1��������PP��h����4I-h?��w��ɜ�W��QiW7D�/8������~�T��H��㜳r��ؓi��F��`���k}0�Z5���r.	���, �B5@Ā���1��m<���	F�L��3�j'�������68O��
�"��{�o�W��i�J�TT:���2�ʘ���223�s��D�� �������G��̬��JDXXUUug��墽4;l#eEH��{${
i*��4�Qc�j��2(�}���jf�'�?jns6�`�.o�Eۗ�3ȫ������V�����{�Ez��1�����cBl&�CF4a�� =�,	ͮ(\��e���YG��͡�.�0G��ݭ���r�� �:��]5����o���gb+�;��L���7A�&ݹ��ʿW!}�j�x	2�;:aҐ"��7��'���Wu���T;�-�ȽO�_	�lL%�a,��FW*4#O5�v���le��f3�#`���~W��.�����s���?t�V	��]�`LŻ�+��R� m���O�l�%"X��؛��¦�; ՟�4�p�.�tv�F�p����)�K��W�Ky�c�k���I�������x�bzh�5�g� ~��m����`�?�E~�а�^�\��ՑV|go�l�>A5�<��#�c��i6<��n$��� ���0�mI�f'�=RO> j�;0.#�褙�G�ytAr�-L�]7��,��[C��0}�A�21,��׋̃�R[uͼ,�O�D��9�6�@��o��+}�H��x�({ܜ��U�f1|�W� s��$A����o�Bery�~��(c�*�a&�ru�0H�8��/�;�|Z�G m��<���Gz�,<%�����/*�'���
l.���L���^���̼+w���w��o���?]�Z'��^�9�=��[��ͷ����h?��~��C����H���xϳ���쌘�g���� �H����B��~�ׄ���7�f�7�$��͝�������5#��^zw��D�7����J2���A��b
�]g�����n�ܯB�bJNV��[��{]֤o9�F�{��Z!�"MMb�d�*�KR�˴=5��OB;k��8z�����[�]����t:�o;�%>��σJͅ���-f�����ۑ���̃MT��|�:�D�#P)�����,�3p����������`��	��2��^������v�9/�:�O�6�v�c�mS�|��w'Ap�ٻ[���f��1������7�RbC4D��5u�Y��~Dϙ�����A�����yʲb�q}
�? Odf���Zq3�>]���݅���{-T�
/=��x���xWo��>�	|�f�Ҩ�9���J�����0:psi_y?����e]�5U����%��]򖋇��ޅ^��e;U�k����:�� ni1Th?������I	
�Z�0�B��d�X�Qx�W�<�:u"��zJ<0�f^�k)nu	"�r���Ei,���_�&A��B�l&p��)���'��/�^����:���.��e�j:���ϳ���vTm���,�:w�Dޕ���qy%�.�����m���D�:�2Y��ƅK���<oy���4�ʮ_�ԛ��HIU=r���ʌ'���Ϳ�����L��x�#�x�i7	�S���&�˖�?�I��C%���{��gG��B�DTlb>VE����?�ə�t��Y�<�����,��==�}��wwT�BF��h�?�S~~��8F���O?}Ԟ�3h�[�5���/3�o�O�Hۈuv�Uon�s�������B�(���Ud�'��Sl�#�E����J��C���P��?���{7rjZ���\o�Ѥ����lh`k�,6a��"�c�k��h���&�o�����]U�W!6Dō��\}\s]�.E� �p�g��x���bn`��S�;��_������!?�Z+y����pv��t�<���٫B�\�+��Qׅ����D�;IU�MV�WOX�m�;��?w>���Ru�0�����,*�;2��~��ŦB�8Ϡ^���I�>γ{{ԣ��9��a=`8U^�d����������6[?p�X�f�dQ��%PeG>E���{2�z亢v�y徲�����j?[��4�y�A��h[Θ,+͈c����ԏ�Wl�.�������X�)d��K���a?��Ro5�"��A\��?j���\\HLn���l~ߧ�Y]����w���射شVV�%e��_W��_���Y�okwTR���=O��־ۼ���������>����Ɣ��ۦ�O�P�$��Z��j�\~NxH�6c�v��B?�W��@�!����yxe�����i��?��b�di&������p��4�q.�)��^��ﬠsAye���-�o������Ud޵�Zہ���	��)��*&4��H����`�eF$þr5{p~wY~�-��+�M�.����r�?	��������\�s[BR������؟.�P^�|�3W���� �E�}��r�����~+�����*'���ҒO��m_�?��N�nԦ�sA�c֦��W@BJ���c�7�t]cs�VI�w���C�Gū�24��U�H%��>~^&���u��,���}�(���\�������Ib��# �-�7��c�z���+�|�Pez��J��H��������� ^�F������?���
�s+���}ί>㏁7�G���J��d���D�g�&*�J�9Ѣ8��c�t=��xK���3:`�&0̴�������L:�_��r�*�.���nT�<�!���n�s��1`Se�����J�SK�R4�?z�"�ǅI����b�<y�9g�`Ҭ���&� x�E,fc��\���ޤ'���f��B&�h$�ҵP����4�#�bY�#�9���&w#FYJF<�cLLL�vI��m��K�=���#\�s�[;��ô[M12��\�����E�.�f�Sֿ@���m'f|Gܜ�c�Ȭ�lD�ᄛ�Iz�>w�C��SK��6��r2z�ޡl��VVRd!�\@���D!�����b�.�	�h6 qLG2D�9xzk�]�Mz���_�C f�ɕ�&�/�'���LMMov�Rds�R� vqs�RZ]��M�Zdx�d�>����`�|}����Q¿l �yJ.�0������ؑ�˃^m��=�^�ӥ&L�z�æ�f��u�d��bI�j�YcD�h�u|�X�{�|G�B�tt�<�3\7g����î�ꮭ��5�PPX(����o�GB�Nj����H�߰�Q�g
��;@�,Z�hB�fL��b�Re"��g��x�%\�;��!�H��{{t]g?�����+�~Um�T2go[�d6V�@o� ��d���9B,�y��i��t67�����'"N~��������>��+�ćJ}W�M�u�D庛<�����h;�|�A?~)��ߘ��Q��:���2���<�ӷ$��GTt��c�\7�)��$�R1(�@�P��ED|�:ْr��D�M�*|32(��`M��̃�&$*{�A����O���_���#n�����`d:�v�7_K\e� �����=�'��\Ć�Hg�Ҙ�?����qq���5�ۂ�L0�C�K�e�kͼ7C�v��q11��0v�c���?8O��0X�ЉY��f����O��c����i�B�I˳3A��4�ɵ��9?�+�Ǿ�\�͓&)l�<	qA�C��Z�l����j�z���{c ²���\}�WOǗ�k,�+�n��vg?�X�
 |Bge���_(�ԛs�{�er���Vh1XH[v	h����,@��\�$گث��QTV�F%wX�P��)&X����P�)1��Ff���iH߱s���R���O�U�&�YD�f>�)fc��l���b�����r��{H\�0!��ͨF���\Gui��r�����еD�@��B��U�R�lR���q��"v���Ւҟ!d�O�T�����C��^�r��{�6\E����M�.u 	��� ��zY9&��X��ǧB�g�����=�IIU֋�H���9�14k�-kxJ&I������q�͍b��x���a�>�����Pm�]����ށ��7�n����P��S��=/O,ۻ��Uڅ���U��ed�\�RVP���+���Vm�|n8mޙ&��ԑ�Q~R����M��B3��_f�<e�^{׮�a���_(d�DK"cM���Kz��}'��l�\�M���p)��j����tYf-9"_��L�z]��B��j�CǪ&�_u�9�q���y^By�,ߕ���VZ���$��g?��џrW�O��{zF��_�2�8��7��[�����5d��=չ��'��PJ�͞���.i�w����EMD��	���/��EE�;�g�i���'�*���}<]�j���� �͘&1������x���=}��i�+{�F�\��1��L:5p|��k�}JZ�>��}w��������k՘�r�9!K�w�4���C\�Z�l�/��3��m�!��+*¬hmm�K1�������\�?�X�/��Q��~	G���r!�'	$���`���?�v���WD1��g�o2����U�|F��@��Vo��S����TS��Dn� w>��T�!��ra��?J�V�,F��X�iS�;�6c`-��H4�H܂��q�`b-E��_��J�Ia?������K:df��L~_J�.v0��>�H�� 2��%9��Jv�Im~>1�z�z̻����N%9�l����b��T�������u��9�!@�7��Pe�c����-�{u�p��=z�z	�^�L�]�ۍQ�x}h�Q�~m�]yN��-&v<<<�J�'�'6�/_J�,x6 �	�"��������.��G�?�`�!�L�����#
V%P��:���N��]&`�74��7!Uh�ȄVue��ȣgc�'��̎��E�l��T�������.�K�d�<H��4�k�Ӊ���C����D�4mֆ��b�;�{�z$q�E���`FQG�W�P14���vܚ�?�ǟ��"�Am0_�.1�v�@���^J��e .2C侥~?���l����)��6Zi�����5Y�`(�6������Z��i{h����w�j���`y�����y���a: R+�ٗp먙o��;W�k��褆K�[F��5����������L����O����3�������rr�d��:1C�����9��b �I�6�oT#в���~����.�\����w�5T�-K�ģlR���P�ЩƂ�6ά_��$��[	3qfy��d?K?	�����-ֻ������gQ�1y�&˦c�i�e'Z����f��>%��i+#赢U�V��_�T��Ts�S^�0e
v����Rf� �6�o�/��L�������'azk��ܖ�<�"�	���O��1�[ؙ�p�6�K ՗��I�#� ����i��Ԩڭ�O��z�~�~D&�L���Xj]�m��5�VY,�W'c��P�;;LEk�8�G,.g*l�6����4hYA�gh��)�M��EԑkȜ�4�!6"i0���^��}�6����R�[U�1����,L �x��c|�J,�
�������edl,�|{y�A���M���X��~���:M'z�V���6�=�mwf)�,~)�]溧mUUr����=b����H@�CN�ό;j��	�gP��*Z?vu�� � S��5Cc�"���@R�U�����[10���X|�	�R �'
x5�`���D{p�~��������Jܻ� ���������XO[��C(Z�ﾁ�H��a�)Wy���Ӌ�!Zh���{ۛ7����wn����xnJ�Qұ����=��8��9��f6�x<y�W6W��k��D �6��6s�,%������2��_>_J|��:�@�	�(��I�V��}�K�"�z8��K�%[� ��Y+��:��;a��ԙ�<�
�3��9��:�[��kL����uvU��e����v��(��)���,�X6�8�maR��ׯ%��Z���>_��q=��4c)"�I�ߍ{J�Bh�ˏ*�&���աI��#�;���/�l)�4�f�q���a�`>�T���s�f�G���q:<2�X�x�V��#�f�X{:�v�/p�Vy���� �Pb���wJ��Z�� ���&X��������;�_t|҄�q�g��:���'[X��$i'�
N��~��:�N��i�'����bmO���)�ܬ+,j%U3;���Y��g7�6��ҭ�z�uבR�?�^}ͬ��خ��Tc��q��.��ָ�Z]_߾��Ml��S���� J�=����B�n���*������|&�N}$�-�=���ż5j3v�pzJd�++Y!�<�r/�ED8gyO�E8s���ԗ����]�eU�O��6�>w0.���ƭI{ �'�����w�[����~��M--�-<L`M��n�� ��<�C����a�(.;�9�jk�u�U����c�`�z�K|�iD茀�Ӎ��k��wu��I��S����0ԥd��i)�����q�$dt�o�0�b�;}��+'R�M���%@�.�YY��3ɹ;��DZ���j�$�4��n�H�y�<>H��ZN)�s��&���4@8;)m{�bp�YG_�X�#U#2T:��*'jfn`_�9TRaH�9O.=��S�虒jb,�ͤ�'�`�,��'~Y;�m a���o�<)�6���TΚ�[��5:��Җ�a7S�K"""�<�<���ɹ�_i<B���Om�.T�.(,Q��Z�@߷��>$��^Li�s%I-ʅ[eHs5���Fۨ:�y`�&�*q�jWp=�T>ބ(�۠��6A�)�i�a^�F,g���Y�������}좊��m|����\u'NQ��Z̖W#�nRn3��Z%�AQBBBq�е�~�ǣ*Sp販'j�lR:�3��j^-�'cl���ۥ-�t�)'��[�U�F9']�^E���oo�'����w�����
����(3���U�aw����<�X�&�N���z�r��=�0U�1I�u�2Y�r��$�;��aqf�W[(��L��s���U�ˮ�ު�X�Z�?є�/l�;��kV\b"��Xb�J�Q-T-��u���$���Sb5��U��V�Uz^��ݜ-�i�������ŏ�31RRR��%��Q�Ԋ8����g��jGEyE�����;Tŀ�Ȗ���t�ȿ������Ww����Xu�'�(�y<y�0������p˺�G��=�Ec �M�'�W%��+��s�Q&+'�Q���%r�j��m!��3,m�Y�j�;~��=�AI�(���"4�쏸[ �c0X�J���l	�0[7��kO-��ץ �����7�#�@t�w����ڴT�YN^�:�J�t\Ϥ��՟-L>��-����X�4U{c:gJ�_?���тMq�y1�����Ɖ��e����������O��6�blIy�v8	i~D�y�դ�|��ж�a��WCJg�׿
qU� ](�/:��}��o�¥oP��f�����bp�HP${����<����N3�1x��j�˛Ǌk��ܗ�g���fK���2>�� �Z(�M���3��n-����Č�j����`ʁ��|K�|[�j��P�n�Hu	��$ƺ&1�#�z<�xf(��#!���'y�S�w��5�#q}+��_p'8pG-��2�l̎UJ�?7��r�[�^���Ț�3��l�#
5)� ��jC%Ϛ�l:�}ijj:겞b�{���ǉA�[�s���RUEŌ��z)�� !n�+ϖ�MG�Sߟ#9F��J;D(����.��.LU
����q���6y�f(��UJ�7�܈QV����~�b�)�+��捰�Z���#�ْ�g��?Ύۺ|�W[�	uy:�=�~[��l�Y��\���ư�&)q�p����g�M� 8�������)��X{�ms��o�e0�8c�r�E�a�H�����(,mV�?�>�HH��3�Vh�͇֗@Zk����E��S/"q���T�����kW�қr��cAQ@�ޞ㧰�}nv ��J����!m������Db�[��|�<�|:4�L��������h��wn[�%*Ė���Փ:�uS �$�q|�?h9��]zh�N��S�G%�+C�%3�)����>?���	�+"=�J�.m�q��y�F�a�k��;�����^?�{��<d��4�x'���}5[�{++|��X�8���}n�#>I�k3�"�4��  "G�nwA����9Q��{�+O��pJ�u��(�2��6�L���o�u�N����y889m�,�g"deh�?�����z|=������Q�qY�0�6J��J$@�aY��߆� �f��)��:��X<)읨2R�R��`�#���§����̓�����vֹ7����<�s;�d�\�p�!�O���pR���tOC��� F*�\�)���fc\ϯ=�cL�*�eA=!�/E˫��v�T����B%*M����Õ��IpiG̿�p�jٸ/:}s~*D�8p��q6�f��/J��e�3K\G�R\�VH��C�^�=�^�pm(vt~p�ۮ�E�gK�X�\ߤ�ء2s��W/Z�,���s�4'K�I(>TC�6�0�������9�6�Q�&��-���{t��F��7�|�_�?����[�z�n������̃��);��n{��������xM���VC���/�����a���=�����Out���AH��u	0(x�H�PM�pN����us��[������"`׃��|��q'���k����q���^��P(��Lk75���ݫx~O����~��ϳ[��U%1�3�9n��2�T��W�+k��wq/}$Q��]�H���h�DN������fv��	D��vhppb�c��^zOOǂ�Ҥ�WS�h͔p'B�e�ޗ���N)��aX�>G��e����k'><�Kj�����|?�U������e�-E��_��5�,�
+h���zs�_�T���a����Y��R�X�|�W	��W�o%���Y��xH~�K��n6oS�r;qx�c��ٰ11}�1t��P��XHH�5s4��uL�\�,�T��O�t�i��]��\��5�e�^m��6��ko�G�A|��.��tx�{{�N��p�>¹����\�NxX9u8��C�m�=��O-�v�"�<�<Ŷ<E���*,�B
���)����sDJa @�9�,��~1���l��|��+Vmr3͖�� 9qr�4q��tg�Þ�^h���X�����d����M9��A.1H�E�eU�����������*�׈A�u�B�Q3�H$�-�p0e��s� _�{�zo�]�}������uXU�k���V���ƭ{�H��Fr��MEbF�Y�����[d:w$���)��PB�!ő�����+o��WUʬ B�Y����8PUYO��ky5Ng�?i��8�����~��f�����������2�L�6�fffX�v5110�ݙ�Twp�kgY񀛭�)eZ���#%*���h��h	)Y��=wݦ�򦩳8-M���a���-�\�s��-��Ln+�BU��m9yz�(�]B��m��ֱ[͛�\��Ȍ}~�N�z����d.��K?B��K��&E��͐ok�a�
�6#�[Kr3�@�{��/?����6A�ynu��<�0�f䃒��v��r�9�ŧ���UM�������z1���,mT�O��#s�J�4�����V˶�j6�ѕ@����q��7<�����f�K�2%C_��밪ss��1���)֒�At�\�>7��@�e0��C7	�U�Y&��Y*H�/9B���B�v�	�-f�4,�:v%V��{����0��8;p~��C�*�T�]�i��@���g�+[~f+������`&ʅN��j�F�*���*���M��[&�����͋IBǔ�p�-Ug"S������w������d�̰K<P�6���E���,}Z�)� ���H�=9�[�ti�(�S��iy�U!�W3s���^L�:Lou��u	�H�T�vT�R�n�9-
h��ʇ�����pFH��~CܢPx�b����)+ҙ�H�ѡ�Q��H���*u�zSXi'7� I2��������3Q�\�,
i��X$�Y�Y�� ��1�Y$˹��B���Hդv�ӂ��-�:"wSs�L<8WTS���&�b/�0'P��/���%i�p$��| o�صXC���@Nq�#�%��J���R|p���3m/��4���e���<F�ߺ~>��U�"m^��+�E9BWg�?�N
���Y�֠���ܕf��}D��G�-g��|iX��8�bL E6A��FN_�m�J�� �{��4?�+��.��s����`!djB91+[h�*|NthߚE��3�P��fK`�h�X����]@�ި�z�O
L��yT��[B�K��&����WU��y��s��������2[��(JNT�N�;�g�ș�A'�rgV�.���ͼN�L�vؔ�G�ݬ���j�k ����)��-X�f-E=a�8����R���]���������\S�@ߢ�#�����<A:���Z[�>�ZI�/�+�u�T���>�OZ���<�r�$����v����3�h��:�+{W�S���	�bS	���r ��I���Ղ��.��첕�k?�w�:�>;��������Iܑ<��S�s���4r8��������|���x1��F��}�Di��L�W���#L���R���4ΰrX%��@*�<Nq,Lv�`�"�7`��Y�_[ѫօ��]نϗ�TRGi��;��o6��H���Y�!r�fMq��k�
�{�U�`�fA�!F��)l.�kaS�":�y�v��m.�||�2���0���-s�� �/�Fߐ�o�-T)Y"�[6ww�y�i6��\&rX�R>I�}֌	��M�>�h�ۀq���d��%���N�˞��ރ����֪�q`R��+E�.	D��q�@F� $�A{�D���q������i��-t�ZU����PPF��E���!o+2)0�-r�R(j6-�ۗ�>n��|���D3��À3:@S�Bq�2\rU�!m�] :55��������EW���ЬL0�E|��v���?6e�*�{������
�9g����=z+�S2%�\t9P�!�:���ou8K&QG��&[*E��:k@*�m�R-�d�f���4�hyt�]����D�TP��z���"y3�b���8�&smmn2󠏾GT_y��A�o��*��@؜�:��x���*�U���:/\sϗR�Oh=�P���mSs��$�tD1��G&����ZY�����_%H�*�B��h)����rC�^[��Ig��ӓx/f�=�XC��$�$(�*r<�pU�����e�QF��KF��W��e���@�����> S�]$tJc��d?2�u��u���|�\$�z�~RP�}/�Vs���
DC�J'�^׋kT����8AN��40�h6�ظ�Q��Zߓ��.�O���<�e���]�	��(�s��@�n\��kaGg<l����f'�u���r�D���b-I���Rf�C�7p"y��n'�~������Q��0�C����a�e��{?�k�4�g��ە��hn:�
�����{��.JA�dp��
�==8O��!ycc�U�/�Ү��q ���2Q|��U��7#�z���R�bql*	w����)�ө�߭���w�������^��?OTY�Rw��;mr��@����}�/5('�V�m�XF� ��l_��{J(6�H�;���Aj ��rRx���>gAM3�0&@Q�!?�D}>& �����s8z�r\f�xc
i�������?� ���<����&���!z��~ޗ�(�!�����~ǂ(K��{	|�����z8#����?0��1���8�]) �;>��(����a�I�@p�w��ưK�<�7C��f�� ���B�L���R8��UؕMܼ�y��!=�W6ujh��[��O��O0܀DUP�
}
!�,�Vm�Q2H�6���-�h�J+H����i6�?"�v���I�_k�J;�ڮ;t�jf�1>2!�c2|��J�y��K��Ιf��Y��)2�ҶA�!��F�*/��s��+A˂��'M���l���~�@�w��<H���qg��v�����F���T�w�#��Nn�x62���gO�׵����BU��Ft�v�m�����H�N�7��'qh�9�Ĭ��������r8��ZQl�u��E���8���0b���|kf��:/5�lđ?�X�(hЙ+y������`���:��|�1�:���א�`0t
D�տd�ʨr�!�D@J�^x�+,h�1�\Dev�W�'2:r��A��ߖ���N��94:88��[��b�Aߣ��x��x�X��ƣE28lE��
����\�]�AF��?��9��.U%�q/��@B�_݉���1�2/`|6�Ȃ�����]az����|	�N���	�W���{zy�N~#�=Y
oO��6��F��Nғg�M[O?���k@Y���ЬC������������|��qV/��4�P��#��(HY']>,^�.�GwkW��yq�#_�Z�GZo�_�\1��%�>_^�Ϧbh�R`^����ܚü&"��?��x*<��c�����vi��#�/����0�LVb�Y1ɚ ]eNNu��K�l
 R����
�Ո�����G�b�/Qa[�z�z�k�]C
g�*k��t�qga��X|��v�]H��" +g�u�����ɱ^2B�s"s��/n�P��m�!��3M�'	�d1��{�q�}�%����P���ԭ{��9�y�d�\Xyꛢ����`0=5'(ٌ�� +0�o��^(�b�Ht-B�o�<R�"K\�L��h�ɀ�|�HM�/�tߪK&��!������i^7.s.�)9ŏ�Q}c��4߬w���F<y�VV�k��O�$��˥���f�D�� �	�
��vX�F����[ϰ�qCDʂ-�J�;/c�Y�c�fJh���Iqw����m$��
*���
F�Y�����b�$�h���&QÇ�N��N�界'�;lIj��0�ӗ$X/_�t9��C��0T� D0f����)���C�f�F�*�{?ࠟ�S[ac����ԯ��2^����Z<÷�-��7��(�~͏�fz��!�A�s�+������p�Q�H#ݟ��Ujk*�Bkm�ry~��U��a���IV	���ң`�ܽ����2a#��V�}� ��~s1���W<5�[��,�@�C%��J���n��#vm�g��8t[�&��n�m�H��H r=�OuG�!1E��Ub�+���1+�l�m�	dp.]�9�-◒�{�M3�i�	�ǻv@�_�w��?�K�5>s�~�<��"�F*Ho;S���<���G���Ur��=�V�N��dK9���O�OC?�0������:�>��<�R���2|5I�����l�����#ۤ��ފ&�˕��x�M�����[���X+"Ф`����Ԁ����}g���0�#�����
<�>��k�k�ʍa�zH�9��I�����OQ��2)��
&��i���3�	,��?�a�� k�Y�C��B��$���d�-pRʓ���.�E��3� ���O��� ��a2:�M�z7e��Ca,�Oo	���d�l�B0�����-��j�.���nT�>i8��VEt=���<���P�I}z�I�_��/.��N�.��u��x�ÔaLR��D=��-��W��pRӱ��e��(;��+��	�`[��� \XB�;����Q��+q�ۿ�q|՟y�W��͆d�&T{5�P"�[)W�;.����&��ʅ�RXFL_�ig�?��@H���[1o�#�������?8���`��GD5�[��ζ��v��6����X-Og^61* E���4)�7��:�]"��_���<�ev]gUJ����U�r@���p��+&H�IB�e����"�O�#��?v�P	���h�O�W#)t*�n���<x��B˕6�؁�>NiW���'w������v	�|�7���"R�~nxd����9���~���)Hh�"?Z�n*��*3�N�j(vb���ټ��t����{�.��F���i�`��HF��|-�b�.��J_6�Az�q�E���ZMڞ.#�Y�vD@��E�_2h�M���?dl��A�Lg{���C����B��-�h����>R8����r]���2/�+H_d{F�n$���@z���a5���0�������X}��̉�5�cp��m���ÿ�[��@��)ֶ�Y�)�G4�{mk
�ޛm�Dh,��Ij�

�JG}�/Q!>��o�����|����!�D4�2����v��|�8s�K�'�C@�O�E�i��@<� dQ1'v!x�$�RknZ�0NS�)�:=T	|͍�`b������}Ľ���ZzI���)Z�F��w�IrXd�]�Z�C��q���A,�cG<��!��{ܣ�*T.����%W	bͦԨ �et �B���r��-�j}�:��c]	높�@·F�o��Q"�d�����{�?��;(���1Tك<N's%G�g�1�#��l���ޣ��^��r���TY�h�/<���KI��2����L5ͷ�����@4,H;Ș�)��z�-Qh���zU�8Z�M�_=u�E��T~�faY1���V��uj�J�[qg��1�@�P�E��9�]Ƞ_|~G��*�v:�X-��Ǚ�P�R�����N�`�˗��,a�'	�\�6q1��|ɸ���C�R������"@�[���K�W������W�GL�f�Kq��O/�~ ��|��U���j��R�?�F�5?��0D&K>}��{g#��������#��@�� ~���LY����(�n�X�N��Ց��c>8�pHJ����dQ8[���e�b�~��0��qe��0f��y#}$��:r�}b�4H`28=<z�_?"�y�����t� s���ӓxq�p�+����&HiR��p�������c��ܛ����s/�l}�����f�Ar��ɼk=�Z��h�V�Ն
֦���0������.Yx�IN7������?�!�c�� ��A�)�-Wgs�\#@ �������������ݸ�@��NC��e ?���w�:�����"����"�sֻ�s�!ƙ����Z�x��<�{5%#�5Df�6�-6��ɾnW)m�޽/Ho=]x�
�҃
ec@$�f�xy<��, �g���p���8�W����<\C�p��L��#�qz�zJ�[�0�U�u�)c���뿃�u���7g���I�6�O Ja�?g*�A�& ܦ�����g�T�z/؄3KА�_F#~w�S�ҥ�����=;�_}��N~o�t1iyx4Q�&;b�|��i."H1V4������pʹ��P@��lQ��ޜ�gM�t޻z荧l���\��ԡ�I"݄U:����1���Ä�GHt�R�7�ܜ�9�n�`��˼�^FQ�kd!b��=K#KxR����?��<Щq��,��d��fPi?�7`�x?�%�NM%�b<:F�-���]F�8��T�yO9$���z��&���n�&�D��v���e}KO���F*��=�2��k4�(4M:��5��Dz��������Hi��.��`��<2b�������6	;����M��YI��r�z�p\���v���/:��nJ+�H�������HV�w"F���[cj�)p[��#*M>y�X�4�����%s�d�	]8b,��{��-��}}Nh�\��������Mƙp�����-���ň>�����·�Q�.��-��E�]cn�'8�"�#�ߧb߳��_Igcb�2��b�E�P/ffE�11ύ����������晩V�\*eæ8W@@0���q"����<ٰ2b�(�!U8� KƩN�Fy����bA�)��n|��ǰf�t�8�g���3�5���
����0�����m{-5T�Glrv�>�&��_��aVT�XH�h�b�Q��N�����Yܹ��b��c�A��@������3O��(T�
+������C�M.�(�2o�T�֎%\����#�k�݋cg�6��;�]�m��:�7�/b,A^��v�˘o��#�{~�lJ�hsN����!T�5[稳�wd^^X?�r�.��E s �rw&�cL�6��	�y��K�		y�����E;1�k��L�cL��gO������^��zQRZRQ�Tr�P�_�Qrtӗ�v�@��6n[�=1ꇒ���n�'�(4�� g�me�n�BMBއ��Ԏ�NB[_��_٤�_�jt��a9���{w��E^������k���-&��N}*�B�l�R��C���pG�_pc#	*���(ǐ�=d <�T+#�s��5Ӯ ���#2�!�������.$�}:N}﮶���~R&�ؗ�x��)�SQ����A\�,�W��z|&���l�4��5�� 2b�F�ܞ,����pOY���֖8c^ӧ�ɓѹdB��ʻ��1�7J��C[I�q|�֘�gc-\cI7��e�|�eY��R�`�����u�ch{|�*?��V�؍�<���E�骃��9�>�mys���F^�S`�=R�t�p.>@B���,�<ڃ�����9?$x�#��0{ٕ�?���ςB�4����LF֦��ѭ�TG�d��ۓ>����w���F�q3��kJ.�e$&v�N+͞���������١�f��Q23��l������D� �A�*(�Nif�o�o��eʣcl�HO&�o�zbI���H"''���j~�vp!���J���*_���W�x��ɓ�,Ջr�������Q��M$�;�Z��ʼ�"&vw�ƈdl�68������A����~ɬ_^�zZ�@�{�CO:(H�coe���.��ª(
(*�te���(�5t�(H7HRҡ(�� 1 ��H�P�yfpw����w}\�׺��<'���9�9Z>����ط'P�hO�{aV��"�ы8�},B��ٓ�B>{*]㊔C"YЪX &�-7"��T�y���Em��1p�N�㞜+~(F�*w##4yڕ� 鵲K&�����S�+ccoq��z_3�/w��<c�-�U���=HUQa��2t��� �א�S��/���o|�8j&G������2��>	{9�,??�P)1��N^&�?�8C��
=�l(iQ��������斍����VV�c%�{No��N��iky�<���� qs7k-*'�ɫf�A>�Q�[���'۠��-�»x8��&ڔ$S$a�\/���Ttx��ۃοǵL���-���*�lܙ���nuZ7�=�uzX��⣚��S���T��|�2j����fo�������-p4uߘw k�/�������E|��j0�s���'ߓ��y,V�6���\o��7���֛^�!7o�{�*_���kr�w쏫�A�G7w�����o~��vn޼��cF�Հ[C����W#�'�?�¶i/�@ޞ@��1P�2��ҧ��./���sY���[������J��?����9*�Nr�Tk	�f�)Jct�������'J �~D�,��g�/�c�f�L����.���s���BM1KΓ�:/p���x�)^� ^b{�ɠ��lT>$�pP�M{�y��Oѽ������ـ��o���$�� ��ވ�Å� lP�z8���&�Q3����H��*$�r�3�&6��5/9lO���Q���{�%tU�h�Y"C ���U�6�\M�����i�t���@V���߽�N�W��S{Mpy1
N��/�钒�v�גb�F���Y�_��_0��/��V��.��ʨ/��y����D���v���k�p;�X^Lm��X8R�����A[��-���TrJ;l����Fי��
��Ӓ	�+F�5��s�]��0Y߿��}�I>ȷ#�O��u�힄�¿X����	��~��M/C����M�ʇ5�ɍ��|�*�r��]�4%?_�E_��[2�p��3��v��89hk���Oá� ��ʶ��$^�E�*;G�8I����2 5{��y"V���a�Q�fn{fw��y%�������G��B�`�2LG/��������ך���e�Z�v����X�J�xO&]���FNשP�fJ��3�������%���qÌz�:,����[]M_�r�6��X��B��ĳ!�н(#��"�yV�d@2Y �񩎳ʥ΂g����&�&$ǭ�z���B�����M
�1�"�� _�e�k6������ߎ���z�^�7
�T�ۓ�o;p�x/a20y�v?3�_�l����͜���6^���{���@��f½>��"�?��ގ�(?��|�/����l�u��f�L$��b�ŵ���$����q���06e%�ld� �����������}�4[��N���S��ЫMg}�ɾW��n�]��/)�M!9�oL�f{�AE��l�z02�݁#���8�����O�H c+� ᑺ`m:B�\�e�F?� Mu�$�]�ɣ���T�9j�y�'3�2ǥZY"��i�k`S�
���� ��6Mx^{~N O�(cp�%r9�Y� �Uź�*:%[������ſ&���ń>������Իwn�^ݰF��CǱY�t;'�!s5�5���
�*��]�ܓl�/�#+���r|]'q<tJX�� ~��J�2��Ւ���|[�F�a�q@E�Β�wc�9���|�����@}Xν�s>Z��3�=)��k ���ƶ^�n0rr:}&��)�� �h��/�*0��?F�ɼ��z'Ɠ�F��nll�׽���E�6n��d;?G&�h��a�Ò��"��2�ۍ��(IsVJ�~�S���_e�*w�|Ww|�v����ER4=��҂��rE�~���ّ��]v�a�|��I�4^;��F����.�V�Xu_�̯�z��^��i�Ͱ�u�ō���J4 vjּ��]7�f�>\33H�ϊ�p�D�t��vh�43�Ȱ�@g>*��`u��L����뗁�Uq�	I��j��܁W���lͳe�,�(�2�0&��g�u�+g�� �~�|����&����A��0R�5��&_��\��JX.�*u)e�Y㦶k12�b�Ŕ����Hl�\֘8f�q�^7TY��@J9I[�k�hfd<[S�5��!]��`I���mTT����Iy��?���S�8*���9-3��!���X��^�f�1=
xr��oI��/{Uˤy�W��C�+�/������w����G�Ye6�2C�a�r�]yCQϷA��l'�$ϼT�Ҿ�\_T�닕X�S��հE��J$������ih�_��	��;��۷���o�{���d�UUq����6��wLw$���srN�O9]�h�>�6��c%�-��ځ�"��H&��&�9_0�crWt��Y)u���� ��2�ÏVL��,�hPX��Sl�W��̄���p���=C�7��_��1�nZVq���Ӱ�ͯ/��/����`0Y�V�.�`�j�d����Nb| �D��]0����@�\�;�I�����W��iғ�i&����u�/��G��:)�� \��Z���o<��d}WG��ܝ����Jy4N�����1A�/u%�7|��>��"���Ɵ�)p��prn���+�i\���X��w���rT�<x1�|��-���jW������9�;�gg����?��E�_�t�g!��D�f��|N������SM��&>�Q<����TmS��9��Y��ۣ=�1��R�,R�Jf(�A��C��bh@-���v'��{��n���:�M�H�0�s��'?��g4�mu�hi|�����F��{����v���n�l�	}����ۆ�2`҃���&�
C�Lb���6Dqs|=�_g�Ϫ,�wn�I+ʐ:��v��OM�o�UO��k2�&��s�?�{����d�J&�&�k��ܛh�禨N4��̎�Dr2p����mp�V�������B�t��&�wM���=1�I�E�8��כ�t[����� �<D�)c�Ppڙ>���0�� ,+8�]���/Ee�ѕ�(��H)�g!�9�e� �q� Ɏ��B�r}�ǅ��%����t��!Tj�z��BT����R	���O5b:~ֻ!��C�����;��^���:m~�K�\�3���-��Ϗ*����j.��I�X+(����8u�� ��r����dg:s�|ɛU=ޭik[��zQ��3 ����\��|cϪ�����Y��u�	aO�����BzgYIq�B�q�ݘ�T�~=��]xUM�\A��&�3�!���A��*��.6J�fS~�OU���&p?��?��`���6��J!��ԸV��k��+���ʻ庬�oT��٧�P��{C�+�c<���W[�����gP�-���/� ��FG�����2g%M�A���rKĞ�84;��0��~v��er��� �,����rMb 7��ȭ3�L�9�MZ��1-�`��
[B>ǃt�JH�.��b,*�˸X���%�2���/��������Ny�8�|v����y��əaY�l "sN��(�� � 9�������	�8�-<���,oB���Թ����l&ϖ�^:���ё����(ȎMw��w1y )�]�ۤ0���vO�v�B���q�*`��sS�b�mmѝ_(�~N��x}4�+	��?�]P}����2 4��T�ТU�����.s�K���C�ځ��񪂣ʴ��a��pQJ݋r��ni�gk�Fgg��L�ͣ�Z�Dy#�������Z���s�ˎ���(�����ݓ-<�a6 �A�c�w�FwO��Y�*�����v��E}+�V8�����e�2Gii4 e�����F�ltG�A�ri����H���8oC���-2N���#��ґ�Υ#Q��X"M�kjp��nvE9�k��o�F-������8�U�����!��T�"-����)�c�R���v�uȧ<��
�s��{�
�9u%%�sWzt�9Y˸�M<�(k�6�i�l�(���Ȑ�����L�SZ�o��X~��D�"�a���8X�ʺ�7�~���������/n�H{�"�ſ�N���9/ؚO
۪�Y�\*c�;�OO��� �Mh��y\���߽i8�pz�l'�>��'�H0mҕ�_s�:��t�0IOb������;ɉ�eRoj�㣏-�ǆ���K+$�n?����+�d���^��%_a��*���h-#��E���ץvG���O�@�a�H�=t���8�]Ü�L�g�AQ"`��RJ��Ʊ���d����&��B�/����O�����qո7,���D���S�A���w��Tsv����s�r�����]���N��*p8;3�����x�ˣ��I�uR�\ҘN���3�^�6q�o�k�ſT=Q��_��?aP\����[
����F@�Qu��8G̎!!Ɋ�׬�bd�+U���j~4с	Wc�|i;��Y��S�~<d�K�� QZ����"���0�̔Cw��4�����SY��*��2��s-B�=��o���BM�zj\���lUA�_7�R�W�NQ��An���m��c����+�������;$Fגb@�	 ��
���s���"o�7/S��ͨ�.>~A�-J �2��?���2ZQk��,����=�a���<�ߥ�N����-c�{��`=m�i�	�[���w/�� �OE�	 \MG/{��r7�/o��f���}���m������wc.ہ�(Y��{�Q�FF?^.��ܶrTp��ebb��P�W�s_⅑y�}�'�Hdd�!j����W� ~#g��ݩG*�?�=�h��˩�r����ş>�}�_�=V)_2�Ҋ\OOc)�p�����oo��ۘ����A���<��5G//;,���!Θh��Ң<�va�����WE��̣$oNjiiAۆ�ڸ�R���{���$k&�=\:r�	7����8<\�ҷ"XEmÜ6@�j�V�0�мx���3R4�I� �z�����f�w�7 �9�Y$�d>_�~
�������RhD7*�#��o�s��Q�)��� ����r{��R����S��:�}镙����mqW�`�l�6;���vA8HF�
뮤�!9.���H`�+]��G3;x�ڳS�Q��(���pn/�[q�e��ޤd>���Jqi*�I]L����L�(q����]lW�������'��A��_LbB|���.ALU� (ћ���j�!�1@'�K��5�BTT�X��������b	�T�*,�i_2}N�nV#�8��N0ɅY���`4���k|n�J>�=����w�\�S��.U[�dK1%9R�jeڡT��|sb�JbӾ/���=Z�����R�f;��eҁ�(�Bd�Ez0��o�,�r��t�Y_8ߊ���wn�
���"Y{��/����
"R�-�Av�6=G���,[7����K�=],������ ���0�5e8.oSy�ק?g4��F)\	�:����6	��;�>�S���W�V���V/���'�HInS ��~�|9JO_���W�)d�?���̓8��X�1A�z��P�8Z_6gQE�N9E3D.3@і���Gٓp�9ts\��$���Y�O���"Ɩa՚l�Fn%%*X~��|�1���{�;�;��n?�,Z�|�W�_��I�j�B�	�v�����+�*-�d*S� F�	��ε�`��w+�m��g���N���c0���em�^ةf�L,����E�.�IT�U&#��f������ў��ש�4b�
��(M�?K��Ą�g�N����͛7�o�q8�J�'f�yN�m�NN_t$Ԅ����M��f����(�<ds��j6���P�2[̔��"D�=oĥe� ��=C����_�����%���A��2����7Eoz}�>HKK����y�MOO#�I~�%�k���[uhM�!u[l0\��_;R��K����&��#Fs��;�!|�߇��v�<:V"�-�"����ڬK9ݭ�E襤���7r_)���d'�_�t��$���*��R<�y�a���������!d��fSㄺ�.DV�+Mm�Ob��<��F��@,�I��xl3{tt��P�4ta��Ȁ[]�++���2C��9v�UL�1#����y�7���K��r�z�����/�K�`m�<]@�@'?���Gf@
�Xm��$���h��(���ț
f�Y���o�ӯ��Yqqq*i��ڥ�Jw�u<��m�DfK%�}���NX�Z>+��y���z���ȃH��+Z����%R	��77'kkk#[[��q`}���$e~]]R��	����"����[�="Ĺp�?;�D�uu� ���뜔Eo����Ï�4�L�s�v������u�ذ [!����9E�C9���@q���\�vz��j
E*�w��GD"eq�W]�gL��o'˒li���"���f?�Ɨ�^~����5׼+V�.�ao�x��"�FP������b�طU�f�s%���(V��i$S4k�����?N���[�^�<׫��˯Xc�l�������oN��q"E�uڷt�|�^3'�@�W�!F/;�I��o��� ��!���.��f����iC-����&��6��:����G�����'�~t��o�E��]e�2wRoD���<Ue�鵘�x��+��V�]�X�g��J�{9��c���$�>G�P	��q.��7�?��u++�,����]��jy�0n�5�VKC�N�l�q�߀;���%�+���c����\g,Ȝ���Ny�y�g��b��(m0��*��2_SBv�?���a=�2�
������+Hi��!��,��-�3��oT�ް�}�iYW��]Wx#������|�H�e��Q%����_��K,�����h������>��9�Z��S��1a�(bbRK���=������L�aO��Fe³���Z���l���ݛ�)n���b=~+�9( �|G��6# �x��w��+e��]����$Χ8v��<�y�������H�TLL2���3����� ���~Kǲj]����������ݞ���>�(��F֣�6���W��Hi#����%�;��rP6��(��1=k�'ȉ�fޝ�Uf;{�@u��^�qM����a���	�I����@k�H����X[�'
؂�|���P�}�9�^�c~��*���Z�`��=��|����ƫ?�}�������u����܆�t�W�Ff������I���&��f9
��-K����0e#�9x���=�{�3�cb�����г��xO=��"�(Cjq�hL�R��+�P��a}6v��S�N*�yg���&uC�	~e)  N���I���#ᶳ�sN�t�e�!�n-��� *7�̈zu�6@�����s�"ʀ�z��P���,`ڀ���z���i�˺�&�xK+�Q͎0�o���'��A�}�@�$�o�0���G�*/dbFzP܀
�5��EE���2�|�z�x�'�%k�Kc�/a-�i{~o�x4�������J�;dpp�pJE��S*�~�r�	�a/����8k�/6l6Ҁ�Af�:E8���ޅ_��_�s�;z2ˍ���5� ��au�B��{@[`&.�y7��"�S����)T��Ǯ���j	'Z&x��L�]0t�A\g��SS�:�.���T:A�	� �%SRO:�<�_⳷�� �{T߈ч7x�#�z��+��������3�&��{u��,������c9�*
L����Au[k��h���G��Ŕ���s��zWW\�t�~�z�ƾ�&l��=Q�+:rr����8���/8�"��ڦՈW[� ೛�7���3J΅|��ώVd��vS����K�t&�u�? ����V~8<uu�u����Xs,W`���9���m`sظ$'�_o�Q"޾�Z<�N�/--ߨ�,g������R��C�x�p�X���f�[q
BD���x�4�ݴ,X�[�ݞ���0;s#�:�X߱A�}��v�^G�U���75����l�����A7Ј?I<&W��
���:����z��(� �c��x�S#Ϧ�Fl�j:�b�<ځ]��u0to�b>�f��!���zns5M|��v�*[���(ɝZ::�?�%׻����xxx�b��C�e�s@)	an�<���\�~��2�~8)���Na!Ҟ\��������h���}��^AE:���R3���4��8_A��萴vr�M�n4(�*��7�ȶkZ�p�$���)�|$r�m$m��%~AFR�Ï\8E�9�]7Y�U���:�џ{��v��
fY������wXXY��`�,U-ՊL���������]��m�\.��#-my���6)1	�Sگ8�l>_bI+ޟjܲ)�����|
�.u3n�ދ����5X=��~��qXFb-b�aʄ	B���mq���6�L��כ���*L�(tc���W�]"w/���?~�$󈧜vƁ�@{�[��6O=��ӻ�|2hSE%E�1�'��"��Ԝ��(��xS�~;����e���Q���x�l{�����Mxv���~D4��\�����_�k��-�S�@�h�i��D��� K�U|������s��Me�s;1���C�i_<yeI��r��>�q���)Jێț^ƻ�~=�N�/��6�}����3q=���[�=�`�!�.��*Ĳē�@'����P=u�s�EV9G��+((���pq�Hz���^�l����)�Y���$o<�]��5f��o�k�;�e�D�;j�S�Km1�m0���[rc��Q���2
�k;�C��^���~Lpg�0�dnn�,��8��H���44Zi��u��U��J����Q{`���Z�p�a�3�]I���`o�n*V�_�"ط�� и�����6Йz�oO �[���=��<�qOy��q�����S_Xh�Y£�H;����H_��j|��_��Ĝ���]YY	�s��A��omP<�!����#0�nQ�v��o���4������!-U�%�������:��}�b�_(7�U�C**h�Â�=���X݌�$����Nd9T%�گ�B"�h��rR�	X�O�ABUC��@'#���� �Kl�`]�v�h����PL�Bm���D����n���OT+�P�C({�����?�A9��upW9�H�2=�䈾G)���{��T�B�� �ł��>Y5n����濟����s��q��|�la�^��A f.���t��t:� ��2���������i�{]q�П(�?�;���ba*����90 �����a����hl���e����3��4�a5`3Ŷ�w�A�QJ��������'a����
`ʱ�+^����W�W=[�����g�

�b聹I��Bgh�C��y6����} ���qɋ'@���WXE������O3�h�F66�a��U�J��5��ܢ����ɒ���QD������L�L�߮;J�:dE�ue�v�5i���;���o�ޖ�b/��߮W�YJ(�=ϯY��tia�>dc�]^���׿w�ji�1�};Y;��VQ�+�^EB��x��D�I_U o��n0���;� {é�OP*R�`�l)Ը�Rc��T���-W:B�pk�ƀ���_@Zk��'�X���vVv��%�WW�Q�[Q��r���`v4ʨ�0ޭ�˔�t�B_�"n{�z��ث�.N�'f�kUc�����
N��֯K��aC���	������4%&&n���)Z�&��N��Ռ��ñ�X�����6��#�\�?���JI1�5�F'��������͍�ܒ����2�.D!�K����E�  �k�f;"�~H���'�kuO�jV�T��ҩ��1�q8?�֘^�ȁq�r����[����a����)�X��+�0�p���<�h �m��{�4�L x�'M^�	[���|��l.|�:�5J�ihb���`-�ӌ9MU��Ý��J ezU) ���|�={���]"��[�|�s7��Z�D��)ݼ�|:܃C;��y�^��^�̋
b�}�X�DY�mE{�sK+���.���=��y��hh�yуҏ�hc��H��ϧ���%���A�u�B��c�.N�m�&͊�	v$��h0דd�DQy�Yy�9��*?��V���?~h::����x�9Xwg۴��Y��Z֣�x,���me%�҉:��E���Warc���Z��9Tr	aOE������w&Ϻ[u���Uc�[�M�rP�r�	�>;�m�2��&�v�7?���$�#��`�_�$�-��V�k4v�X!&�Q�CI�kT����1�%V6���-�(`������ۆFG�Pj�f�	���]�b���âu��>m �{8t�/�3�?'��CŤ p��yг����s_(y�٨R��l��	!]�#�]|}j�����\�{��Xm', G�=�6|��н:��LEђ��EH�`Y<�B���R"Wr�\R���v�K��	@p6 i��3��(�ͽ�>v��0^�3g�,��ѣ �U��ʣ���kk��n�_�F��=~A?V�A�C����uG��p�AS8��;��<Q�f�<�<�P��Z�$~:�<N:-���O{b���zP�K������X���������y����	Rń�
�)�aQ���
�����޽{ ��i�x4��u#�|���g��@R��\���?��o?�^	�&��4�Z�-��ݕ&��q�p�<��Þ�_}��{��7uri�S�>n{����� ���6���D�1V֫�yZ��_� I��Y_� ��ge�Jd��Y�U���X��Į�����Z�X�_���l���?�"9�� �M�w�����O�PN`��'�������T���H��J8iW�P��ԉ�^��4��E������4x{No�	�)~�^�^���� %W7H9l�SbV�J�{?�|�I�Cj/E��{Ɓ"ST����h��D���zR~Iɰ��ڥ��%H��N� ��e|P����%�<��5J�á�&�*mb.q<0�KO��&X��׸�+�$y{{���ߓ�$I.�c��|����@]9���P�Z�Jc��%��K�}�c����>uD_9c���
�J�S~ު1���4�<8�E�v�嵦β ��S�2d�j�� e�d�d�yG�
ٱ�bX���W�g.�F'/j���g>�ty��-�E�~
�o7#����
 �AT�(�@x\��	�S~zz�{�_fS�pCE��Tzf�=h;$��OfųM1f_uѷ�v�7E����� @���xE:��Vx`ǚ����� u23/il�ߙ�
��X��#���Z~�4�4tt��i �GFX��4~2<����Y���Z���߅�^W;�6�.���v~�Gκ�-\SasM��Q�8W(�ĝq�KxC·'�Z��,��~-�gs��,.�\ۻ{hk��q�O�)H��%x�[9�(P�Lm��e����mݑ�T��j��ʄ<Kr��V�u�f*
]޸rV<g����M擛�98�ʣ���YO�٩�u� 1I�#��­TW̣cc�B?��\�*,޶��^nַs<��J�a��3��)d叽�����R՞I��S��㩥�{�2������ԣ�����!H�n����Qe v�OII�n{�`�ܨ`V�iG	�@)ł�M4�͓�������-s���tU����L�0>�ݱ�Εm��x))�����ڙH袠dwyq�k�r�й�[���L�@{u1���mu'I�229�lu���i��D��JY��}��#n�#�N�� 뢾�M;�HG5����E_����~�����Ai,|YJ+B}>�c{����[,|>/bf�O����$=�VP|"�zl��`cﻵu���3��}?�����_�ġ�b2�x���sth�E�\����8~v��$��GB��8T�!�5�e���E6��h����&cɃ��J�M�.�X#o�M��c��5�.V�q~��5��n���|0h��T�n��Lm\Ȝ��2z��F�gt	#����Y��1��8t�����o���k�/�`WV�&W�?>?m^5��� ��z�d���C`>Y3�9��*�W�id���9:�ߋ�����į�����6V�V�+e�M!9�5jt���X����9�?�Ф�����#�ư��7�(	�|��C��xmF�]�ӝ�.�JO71���lMF	2�����T<0nq��U��v�1c�ފ.W߃�����Om��o�Cᡫ֒\��5��VCe� zoYsss�|�+����-��䁻8��4�י�#I�t������z����|�����7���s�e ��Γ'㩱>^�y����C�^E�R���|��C��;�]�i��n�=&e#��HUGǊ�$�x/���㼹�9���e��PW�ω9�9>�ӚG����^����Ο���WĔ�?l����سtgɊ�F_��5�"��L�2��C�ۄ��;�d���Ӄj��Oҿ�bMP\̑�σ�����������v ���Lj�El���4�g� ]d
$d�F������2�K�1L��K�-_��� ����0�3�Nߵ�.�mZ��4�d�\�D>���u����$��xhZ�9�Yİ�+�>����{�NVtT�#I`�������#5���;�ѵ/��ĤY��W9�wV���j�-B1��CQ_��� o�=�s�_C�[�Lt)�Z�4��~����[(5����l� |�Pc:�q���V�apHǸ(�`#'v�9"NF	��u���`�R�N� �:g�E��ho%�����ŷ��z��b��So4�q��IJzM�K��ߦx'W�溱z�����w~��>�����'����d����y�(�~Iy�'��O�]�#5���D�%�{���%A���m~�İ�W{�\����l���A'�tC�0�Io�����0���Ϳ �#6�t
23[T��[Kcn(%����>D���r�p�"��+�2RZ���������!]����7ϟ��@E�q: /���)�?MN^a�q~i�b�R�eveR�kZ��p��8��n5�$O^$�u\V�F�:��d�J
������������뼵[��-���Zͬs�_����|��"G�D}rS����ޱQ�9u��G�����ӠZL���*��|�F��4T뉖��ؖF�����(�
������r�#v�с����LPm7?'�A�ؼ��K��l�>b.��b\���Z�,��� �Ed�v�E@��k�j�LK�fư|��+��E�B,m^��8,��»��j1
JU�;�zj�7�0?��lJ44�)�Y�p��>\V����s�?����u�9T�1�΅*�PlaY4�(T&t$�$��
�^��i�&T���S&RAס^t�^|lo	Uu�^��S�ӊz �!e=7g�R#y����p����7!-EI,��Xq$���Di�'�Y�L���6,7[4cטF w�bXf�å��ӏ�+d�u��;��䰸���'��U�<>����h�):+޵G ����E88�q�� �,��{�Ms�;)�����N��[�C�U9`�{{�Q<�dO�>�^���X�h�OG�VE�H�L�n(�"�,QEq\�z5⩊��~�uu}�V;��1ӹ��A@u���~�����V��}mʠ�zê�ZUk�ݍUjs���]
n�k�75�mU���vě����ĉi���9dco/ #c��AK`�́X�+(���7�q���lv\b�S������܊�A�kV(�@$9�O8m,�5��ݏ�$�����+�+�l/�'J͌���^?]���v�sc��Y�i]� $�)�ݸ	!s�P4�nx)[j�Do��.ه�>\����&P�v�I��K��*�Ҍ�e��e�B0hog��\����L�ih $T��\���y��VJ�q���\�Z,�@��G�x��㣳@��o�F��=06��W�Dr=u�n���6{�bbرf�,ZIac[j�2�������ht��3iQ����� #��W�6��5�u7{8�E����V�7t&�9�mʷ5ǿ�<Q�����]��iLܣ{u��ٳP]T[A!�o4H��� ��Ĳ�ƀ�;������j�t ��3~A[M-�P^f��S �5�>�w�}I�LN�=���P����fck�;�a��q^Hl���>�]���F�`f��|��F8��l���/J���]ۇ�֦�z(���۾�|G4}��BWn��S� ��J51U$f�^��ɇ�����5�|����Y���A
��e$��C�w.Ć\(�&p��L5�ڛ;y��}������,U�/�b93�Qt�8�<H��M.,�� 7����$��S�ZD�NY�O֮���lTgo���D8�$�&�p�ʦ��]?��<�D�#=��UI��`:������F �7��
��<
��x���[UME�Е��2�z���ϟ�⃙ 3��%D�U:
�O��!I��/fgg�k��Jj���������PI��ڏx�i�ڑc=�ު����d��v�B����,$����O����0+�۬,����7��v������{�I�Ц�P�|RX� c��V~���Y�*�3@v�;��2։�"���а�E�XS�	��NBe�Z\���G�E���S���e@�&n8	d�m����������xXa0]_��֖�p��^�K6�%��k��t�"y�N[wߏi���W�{����:j[�L�x�QH���<z#�?E�*�I4��`��q�ߠ�e���}������15��E�g���U�I��nwI�nC�Zӊ#v����{�ɡqzM�OV�;\G�@���*,��QjW���z������(��v)[`��ٵ���t�w �דz���;�M*rkR	ijB�c�Fc}�O�P��0��S��&D(�bf�߼gn��g��W7n��m!����j����D~c����%Q���@�R�|y�t��=ty��{�z4��0$� ����y��(㬹ߜ&���OC3�8��ǝ! WP�����T&q���"��_�� �.��ģ���]#�nH1��v���g����!�@�d	�Bz����$!G�ׯ����':��!qxR��:���)U??q�ۤ��Y~VJ^��bN�����ySq=Q��>�Q�e�2ν)����vpȜUWA�"��u����"�j��]8�;1�Yekn��{W��Z8h�i���! S��kvD�^P�+:�t��F�g$���H2 �:�Dݡ�%t��Ǹs�:�����n�m�GAqq/�Իh[Ԙ���P�C�	d?�K��H$J��PH�"�o�79��]�K�:N?hO�`�S�pPS�N?\�h�]}�^�Xz�����F�v�pO�5��+�l��Y�+��Ȟ��6d4߁]�G�hj�%�9D���][g�z�T����ד�,�̝���ͽ5,��,�ږ-c� _n��Elj>V���P����tu��/��s�HE���=��---
]���HZ��75���.0B�FFŀ�A����������}�~��2���|�}�*�q�)\���}�-��[	 ]K3h�{�����p���ܓ�/Y�+EzVTw����ј�h�T��z� f?M��C���o�.�ņu� !c
��c�GF�0�{w��
��L�L�
-��a~����
���3 ��!W��Ư&aU̙���!l�������M#1a�LF$+v��S�LnE7!!r��J|�V8�e93B/nG~:���P?6N+��U��%0�?�ajCF9��^���y���\�����[
7�O�D$��ȭt������@�҅��C����ᢪ	��F4�_	�9&;++YNNN�i���F	 ����e�� �n�8a1_!af�Rq>�S�R�<���Lx�f��0�5�b���e���B��7�2xɭ��Bwe*�_fMϮ#�U���ʟ�&(��e0��9>9kJՠ.�YE�x.''��ߥ׏�C�uE��SP��Y2jt�~�S(6U7�J��������THv�R��S|��4P/^�nN�Ra.���%��Y�������ʟϋ������֟���88����7�{/ 9�h�m����k�m�o��+�r`����re��5�S����c&?�������Z-����%�=����ȼ>�����/��^���zhh�Âo?b���}��I9u�˃�~��;. �?�'����A}%�b�xJ��+��#ԡ9�I��ݴ)go��d����'��<��P�㥦Y� ~�Dv�{A�G#����Vڵ��y��ݷ]}%_~����l�GpzbK����x�1`�.݅�K� ������֏�L�1h�<�Z���#�x�r�;���l7�WN�.Yz{_9��m�%�2��Pű�[6{}�#*/S��2A�r��X��w�^�-������ȉĿ�:Y	�e	����i��^K�~�۷�l��U���$����:oa�f�
m���R��qR�Ƞf �ݥ���0��|�ug'���'�Β]w�^��.���0����Ǎ� � %C�b�<�{�8m��w)�@�`Re�L������Tg�l�E��&��#�Щ/U�&<`�X#̾5لڅ>�z�j�4Yd�2�N�|6���crXhߺˣ`%��d&'t����.A��5$޷mq��"�/t�!sv��]���i�JWI/5{A��-�⫛�� �۴������������5��0	h��20;�cş�%���k����P�+��h��v7]o~ɍl�c�a��	ǀ4?���5����4��� /�b�6�7���lP����nM`��p;X
o�x�7ܕ����f�����K�n;,l�m<(7؝}7�)YuDZ���ɽ4��e���RdZr��(b[G�8�̈��OE�O�����t%�5��#���c�H@PP�����\;�v�T���ں]��}FX�
��������z>��.A�q^(�y��.�&���7#Y+2���}���Y_�c��r�Jtg��_�\��ߠlo�Mv�����Q�G����/���?mFI�Q�8��=�FH8𝛇GR�����B�|�S���q���á����}l�c����Vb��B�^�\������̭x<�`��g��͑�Ӛ7�A��Hp�!BI3~,E�ѻ*������� ��@�m��=}\�����H�- �'S`���� k��S�^X�.1,����;]����MT��=:�*�=���5�E��.7Ut���.r�XS'�ݍWS��i�E��d����u�T��-��0����{��h�݄-��&�tgi�O�T�ƣOa�P�/{�N<�M��A]���-*�A��	LM�����j0B��
x,�Αdu�zQ��*z��γ�׻q��o��
o,�{k~0�ڸ"�~�w�+�jdz�j40��/:��*}�V?�֞���D���Ȥڽ=r�GrK+�m��91v�G10��������I 7�/?��l{y S
���:hqU'����'є,#^���c�̩g�_�����*^�.*�4��7K�NDA����l�$�k�lq��E@�=�H�(_� g����t����c����h <��4 sZO1z@�	a��EEE��W�**+���Q=��80,�������)�R����n�����,k��T���>-�	%[��G2���Y8����r��<7H��b���5�U��)�k���i���OyHmF��+@Dˮyݜ�Y�����uh��R#��Znnlć=�[�04��wV�����t:Di�[���������<K�?�w>�9��9����5>�A��c�̳����G�Np���p&o�c��_��]�p���	h�wT��\�ؿ&>�ŅQ�_�#@=��KwPEf��r���X�!Y�UQF8�%��=���9����ٶ����N6�=���W_��*�?�	%$�YRD��Ai�X�DB�S�A�C���i��]����"~��^?�����Μ9�yΜy�Wgp���s�Z�}G=��NMv��)��K�J��8J\gt����w/)�o@��g�q��cD�7�&����}e�2�`��W�VHF����Y���k_�?/ѫ�c"V��6������Oę�PR�����,'x��t8e�Q׻��G0�ȫ=d�s�bmOً`JO=0��y�V��oB��=,)�E)Hq�z�IҫH.��d�m�,��hfkcm�}�5��~5!+�����9R���WT� ^��φ���P�����&���	55d�R��tX� E<�|M�����
�w��Ԟ�|z�Ĭ���'"����$�}��뎞�#W�yπ?2��k��������'�ɷ����l]�'Ǆ>S��.�;U$��帉"Sv��VG�|��2�vh�w��ߦ�8��L��w��~�Gt���TW��)����u��++G\Ü��	�@�Q�*�U���;�,=���ja+X�Q�(�(��H�ȹ'�b<����1��'�������D���?�-�T�x9�k'��҄���}i�~Af/C��׶��n�6���Ю�F�y�d��㦔Wb���QW-G�Hs�g�i����<:�Dz���Hs�b���M�Ν��;F���
%2WM��Kݦ T\s�4�$��JZ�~O�Ù��k��5T�ʁ�©�DL�`Cd:W�cc�z�4�2m�t�i˄`/ ��tu��q@g�����<�H�U~����l�x����\5 ��M=#�Nv��,�*`ד���/3)��:zId�z/��i��~}�w,������6%�'����w�1���is��$�uz��.�/P<�ƱLw~��(;;�	�:�v����<�0J�*y|k�\5q��҂l���ד�21�`�K33�mJ�Q��i,%��O�k�-�&��Qrp��ay1$�;���u�/
�gy�M?͇DҦMq����{�!]���[r�3�<��$-\r�*�����pnJ[�`D�Щǥ~����x���{��̓�������h����GR��kv-8�@n�2)�4��uϰO���T��Ȉk�|�S ��'2��O��XܾE!Y;^Kn$����I��f������PWq��M�(萬�� ��ëÊL�����]o��׵rx�l�kc���Hx��m/M^~��M"��w��"����h�Mk���g��N�3�^�Kx�*fR�q�YX�Y�gΝ$틝+{v�~6����� �sC��cWAbx �	tQ��V�p'N�W���ٛ��P4��+l?�(6���n�z�6'5 ��^�]��i-�6�g6�უ��j.8^���\*#>��Ǟ��2�Nֺ�g�m#V����\���ù'���=~��^bXR���a��3_/,(�q�E���'dfV(�ߣH����b7���0�rƈTy{H��B�C�Q.ͼ.P��Sذ�����i��<kn��� VOU�5kt}�U�"J��z�`�\C��а6���eۇ��#���Z��y��,`�-�ef��w1��y����7D�r��o�mt6� Lr���<�s}{�?�3��A���]�i'�fӲ-J"ojWW���҂Z��;��� �`���NJ{k����d�?���Q�XIOBJ��ɞ�K�6(���b��n����[�#,���:�--6�5q�2@�f�jD(��tMhyu���M���� �d�}���*o<�
Xcf�E�L�B��,��������}���#��O>�C
�v:|�g۷�E�� J"\꿧Ֆq��ui�kx�J���5?e��p�;���Qr���-�	���k���+���^Ű��g�F�V�ԧ���)��(9���$`���؆J�L��s�ز'�H568iz�5�{)��̺{������8�����á	���)O�QY�9��6ؕ�`�4[y8�ΒDy3�o%�.��.ץo�b]�^V8��3�:���X�x��V��=�_�|T��xg�WflSě�=�xRte�,��c�o^~�Ggr���X�UJ��}i�;�R��� �N��E"���&h�T�%˩�-�8t���d~�/�`P�r�'%�M,���S��-����B�d��=���az�7������K��]Ǝ�8�f�vP�%.�;$��֜��?W���k���u&˩;扟m�b�&��Z�|^���aeeb��M���4���5�k�`v7R�7<�0._�de����2Q��8
��e�ŭ�6�V	] ��n���B�3*ؾ@{��n(8vcT�B}=�ۯ�x�����˂C��v�5nypK��#l����R�\^yGB��mʻ��^�o�#�؜W�}��掆:Лݕ��Z���[����(4�O��F8�Ngtj�8B�bn��2��Z�xM@���� ��3�t�,H%'^{���駗������mm�S���4�ͪ��F_�?wl�j����ޑ5c�0��O�7g�_��u�<�]7Z��;��bз�b������VC�O�����.�������0Ei�5}���t��w7���|�qά*����ő���+�<�~A<e=l5Z��^����K���^��g�r��b�9�M��g�
����}pbPߟ�?%j�Os<�
�(��L�di��E���3��؏�Bஓ��l�T�,F}2a���!�_���/�ȫ�R]ΒC���N6%a��G�����I
���w�XHC��� *;"�:;�i>����+6�ʻq�:`�9]Դ�=4އM���j������'sU-!]ָ�f���K��5���Qؽ���@������!0�C5f�m��ڦ�Z�C��SS��o�ѝ�(�����+�Hkf����	��)���x��^�6���nd&}/�������I��I���pv��V`r?�aJT�0�����W{;�-�;�c��
���q��'��<�rO�e�rUMH�'kr�T���^�%����Ǐ��Q��A�.�?�Q���Յ���gs��ܕ6
��H�KP�c�:n͜X�͉����x�����Z�f���Lja����9�����o����sF����=خ��Jy�e׹<?,������ő�A�1F��џ�����~[ݦ0��C�D ��6Lc��#��X����j1r� !1�Wo@邏����ݚ�y]��/Vŕ[9v���dӥͨK�ww	�����U~�I1�P����j��7�Q�x�S:�̐�7�r!����'ۤ����n�ov��	��*&7�T�d��2#����{�Ħ���nX2��0CI�R}0ť�k�O+�Z��,L����V�%�;�R��-���SL3эv&���R�V��J���(��:�w<��E킻m,�y��-���Z��C�7'��s��p㏵���>Ϣ�9X��d	�0�)��&�
M񮷱�ǒ�I@ۑX�KXԌ`BeJ�����.^�Ձ.rO���L��,�}%k3vύ��+��Ϧ7�w��OT��P4�I�.5������>4�2��Sڤ��[l�:<K����uK�kc�Y;n�u{R\���md݅Gs1sb�d,�6l	��:��U�{��
5�תTT!�'���,�m���B����5��-�C!u�/��=���4�����mK�_�<.�*M���f��.`�iƱ��K-#*����y��3LN����~���9&n�X�9J������O5���E��4>��By6\��N �r���SѢLq_��]cl`w��Vz##{�����	'�=�a��;���]{���#V�TA�,�W���1���L^	E�K'���0��`:��.�:P�ۧ�P�~,s���\�b�~�w:o����-���q��w0�^H���s�^~��:jb�^�?
�h���V��0c�lBccF���g����柜S�w���&l��z�(��g]���8�T��i=5�O���V��zs�?�t6/��Ll��<�'3����A8�<j�k<�d�ږV��u�l�.�4tV�(Z'̎I�_��>�8������,��K��vv.8!nu-970��eom��e� \L�$nP*r��(�`9i��i�q|y���N�����Z��u���'/	r �;jT4�R���i�K��G Ŧ��o�R,�Y���
�G��"�nb����N��o�̓�i�,+����>�Y2�Y�6	�)�u'X��@	w�� trp(^
aX��c������u�Z~�L��ҭ�t@������;�n�yiDl��l��6
���}� Bu��(ؾfS�c2�~E@������:�#��kyq�`qK-l�_P���������3��<r���Y::�~�o�p�kQ?
�<�S��<����W��wF���|�B�7[�:���1���!��#[�0|-�\�kv$EL˥99�&
���CT�j4�)B��+���7��^u���#C�3���6Y���R�e.ڟ�l���d��>�ĺ� 
����Y�(`����J��ݞH������:�Ɇ>�D�2w"�VEf��R��ѫWG�'�8&?�B�.=>v:���ȑ�i��ƻ�Z�S����v��m�c4����N��{�<S����N��y*?�9�G86�`ѻ �B ^Ƿ�@5Ns�5~h��V���=	�*|�O�Ǔ�w�(�z|@�Ǜ�rP��[{e�88�B	��s�0
�{���Z8Q�Q��$V7U�N,0.(��}�v'_���d�ϲ-g������kj�-��g��������}�.�V�\����bN.s%�Ae��)�F:���%�m5fkKo�'Hu�{�~1zZOU;vL�A��Y��p�|�P��fs%����Ǽ�|x�נ�Noo���Wh�������S�8�j�|��00�	xy
�'*�g��Iw����	���@�����ox��uQ�1�ۇRL���cP�����zܳē�5ν*@���� �.v+'2�/����.�)*�vh����Ǿ�j��d������_�ƫ	$��p�e�V���.�a��rP>�T4�ш*����!"���|��F}ҝ�Zş�������^��RXq}��R�zE"<�Ok�/��f=��⮗�������#��X�M㧺zn̜�h�U��c3kȠ�*R��x��Pt�$N�����/ⶌ��]�ё�[�I69T�nc_�p͉y��	Ji�ȋ��_�0�>W4�ւ�u.@G�`��4�3�E�r�3Q�T-v��'�%�g`��ݮaN���6����+�#�c]Z�Z!9�&��@X�bHhi��$K��}{E��U�B����6)���.��>����n^�s����k�����R�D�c�7��&j���D
N�����^VC�:�
�F��O��^�8�X��]%�0�I��n����w�ݓ�p�Q����
*�b�4�[���Ӝ��YSD�'��+Z��kQ��*��R�y�" �����
"Ï�{&�W��湄��V�.�@����	R"TK�zb���QP����7�� �^��j�G���Z�LG��Qou~����߉h�">�I���C��/�w��*������� $tO�]�P��^��<%��� egHć�É���}c��<�(:��#�R�}D(���HA���ø�_�~���3P귦�XR��g�{��Y����������-�*C�w��"	K���T�ˉ�� �>!��N\���f��3��s~.�-~�(a}�"��ܚ��^B���<��		���)��r�����~��Þ�~ s�� 8j�	Q���;v�6��"���y�zOzWl�-���&��]��>��1D�[$6�܌JR�<`+s��<[)�W�G�\C4����;ܫxe*{��fl���%H��;|���A4~&���,li�qC��ظ�n���tje2vf樾8�a������ɡ?F��|W�kȓ���h��6�ũ;&�	�H���~���Vj��k}=z�y��/ʷ�2}�J�'t��	Ҟ{ T�0����>0��M��|�G�~�~�mP�-k���g+C��BƫR�ǧmyy]�o�{��m�Qeh�z��Oa���V��jxP����r�Z;������ܕ���OEo�uqWS@�3�A{�H����8sFs)Om$�/��aT�;/o�������c�#����JL��c����P	��ZsqeI����Ζ�Aa����b�w���(��=�D1!أd
ʇ&�-��/r�k+�[<��G��TM�n��zG�Z#p��+A�6n-ѫ%������Ye����<C��T)���w��E{�� ɓ��� �Iu���É�XV����J��l�٬���Kq���/��E���]	t�('c��7�kbYY5@Լ|劢�`���܎���î����Ù��iaiJiB��Qv><���wG�Lc@�0s�t�%Aۃ� ���/���Er]"u˘��]��}�S��U��V:y��g�w
-'�ߗ�R`l�om�ޡ��8���F���Rt����)L}�+HLCU5
��ad4��J
���?d3tLș���#�f(���k�N���أ���>W�12\١���3��O�g���qU��<�]7t�\�H_�J���U���z���t����G߇=x w#��H�6O���+L���m=<���o߳rU�>R^~����nM�u3n)h4ZA��5�9�*���&�m��]�腕'���h�Ј��C^aᒑ5������li��;	�6�;�9Ɖd`����)�s5oY��q׮�}PN�M�z*�!�E�Of9����N�:
+�����L�-����=� 8Ȅjk.K- ����r�󊒲������h�-G���6KY��O�~�U~iV�C�?�B�Gg�[K��W����S��,J|��ɑ��i��\�o�B��{'=nyyy�LSUُNp��3!L��/fc���a��n�Xm��ɋ0V)�8.�XX�s�)�^W�tI�q��ɸ]}43K���G��aBhhF�n������b��R�wC���c?��񂢢e�-"�]X���|�Qt3��8��F�n��{�<s���f�s>�l'H��>f���ي���Qܽ�M�vV�rg<�I$�֝HZ��p������b��a,qrޤ�x{�o\7��ɍ�8�ʠ�zX��V����@���g��_ۻkB+LC�}��|��� s�Y�5[����lvCL��R�wY�����o��������$v %I��ξ��.G?:\h=rFID#Z��	����5���h�"ǎ�f�:(|��w�����Lpf���-}ym����\��`I	ｵGT�z���[ʗEm����pd��[��[�X�c���ǿ�w��������5��&�^�NY�SR�n\:���>%W����^t�w�(+5}��13#�(tFݪe�;��u��p���sؔH��KqCXņլPW�"��.EÏ�����?�%Ɩ}�l�����*�R�Oxdf��'��"��>K,���|<�.�|Lom=�
�
q�>���{(��7>���Ւ�m�(@9�v�Ѷ�.\�O2�u�/}���p*��垞�V�N���Y����/�O��ygy�z\3^�f\�_�G�O4e\�t�n�3�j8h��C#M���;�̥D�NR�A�6���YJ<^���|�	gTE|vS,�E��.��$���m3���~e��W��/m%���c~�VlCH'�� ���6�t����Bŗ�$aVy�阯9|�%P8�������B��1Y^����rD�T��FN�
�����.�ܷ���1�mz��I'>&��<�5�t�\��`�ݗܬWՓm+�f��+Ԛ!4�7�W��s�챠5��o� 4��]�`���-~�n\�ck��dm��Jt�j0��HEl��a���0gݶA��_Wf�0������u�������X��b�2:^�~~��h#�^�x1D��L�&�����C�PX���b3j���A�ռ��Pw�aig�z!L�06�Z��r�5i���)2sJT�����ntF�����C��ABy��bܖI�<_���<�zM߳C�c��E8b��i�:$�!y�Dv��[���+�6ϖ��t��ᦄ���Y��'XE�aS��o�M���f��� Cfk�w�K���jb���WQ����X���܉pqM�_���y�@Xm��
���H��{�$��x�N`lF,S�z�=���/lmG�S�>_H�TU�_>n��z���I~Dp%�.a6GKm��5��m��HɆ_���K�o��P��>11"r�e�s%"9I��t�i������&�ΰ%�a&-͖�%k�m�ǎ������Y��/ x=��႘�='a���Ld���\���EȺ7"P����"���?�=��=��-:�Kg�^��6���9^���m2F�o��P8��\�+';XtI�Û��^��:�Yg��%���M�j�m�g���8�I	6���9X���s�2N��o�B�Q�����ņ���m*���覾�HHI��et��ɍHs��>�suB����vRc3�n�;f_�#��͔\«�jkD�ˊ�������V<E�06�.�$B:)��F}~�3�4E����P�b�;#cc�K8�h�tS�@Y�(����-�,7���jg�t����N"�9I�׷�7���z��b�S5\�ss�a��ϼim�q��bB�K��\n���.�fU��O�U��s4q�bk�,}�� .֞P���L�˯[�:�e�8�m���Vz�ڣ=�F���qA�?h���7~���iC��W��O�B5����R�*���S����`��NNN��ЛU���x�f��l�� ߤ%�	zH��z�ߧy��p���M�j!֢?1sm�L��'*q�{EO��f)n��x��S9?��C�S��3�z��Fw0oZz��.�(�W��i	x��s��=k��i��basG��q "M9��Tۄ�%'S��U,�ޅmz@����k���cd+++!������r��pg��U�T8�_��B"�p�'�q�O���iٛ���`kr���$�I�0�	>{5���yG����nN\��/�3O�k��}@��D[��\=��V��S�G)Vr�Y�����C��'�[� �O�J�Btnmo�<�]�V��N$jiO�>�w�S1�3�q�Z��Ҵ��quY�:�K�zl�����{sAK��˼#7��9s23O�9h�F��ϵ��ׂѢ�P���7ta�7q�o3�N�3������{��ш�΋����FX੣k��)����M�ou��E�S/�F)��A"K�
-Ặ|)��IC�`|j��,���Bֵ�A�W��d�b-�W� AĖ_�M��>s.��RF�`9�Z��,L���ԯ�h��z�r�=Tkn7�:�fz+�6X��������4�'z��8�A�y����R�������ZҟN''�� �*<$��#rn��*����Z���(�<�H�l�iC�9�J����Ӹ���u������3�13�4>=�y�q��5)�^��Ɋ?X�!��0HV�>����/��gff�R|��K�M&�ʃ��\]G�L)ޣ�i�=,	�=�2=��J���0!��p\�W^؞�V��Gv"0[8q��`^@��L-�#���.�@�_��'�����\e�2]H�a�O����h���4���]��څdK�:�T^��ƍ�vḷCB�/2�E�-��i���y�ڛ;-*��p1{����455��J���>j���`��~�*$����Q��P����K8cw�JY#[0B�K���o�fjj��y�<��P-^�1���f��$'��^&ك�!��V�G���8�GGW����o���� %��-9��oO�a�"�8��|��+��~�
?��@2ZV����b����]��Ǜ�K+]_�XX�>����L�އ��^�*]��Hf�����GvrQ2���T1�$dd}�u~����/�s�=��Z@Vp�%.#��l��T��=8����FIB�p�{��f*T;�Y�r{�F���ж֔c7i�2��[�̈́R.&�i)Vƚ^�~~0.�\P��|��?o����"�ǧOuс�z�2	|[>tpS����:���0/O��y+$k8�*�˷o���-�$t�s{���A�7�B�[�=ys ���r;��p�����]t�l���D���AK�ї�M�hƪ�܀6JEZ:(9%z[�?����n�Zؚb���D>��塳y �ڮŦ8!��p���\���I+P��h[���>�8�`3�q�W�aդ$��͖�	}ʜ����=����o�)4����_��g����\ޝv�^ꍃ����F�i��+���I�^��C}��
�l�xxV�+^���|Ms$Nf��;t�0�Y��=ٞZ���;/8/�q�4��s��B��Ѕ�<��&��G���џmMCC�񵍍��b��,���Sر"������nk�3}�t�.zh��4(N;������]\�=�$���ƥ��M���6ڊ��\�j��{Ez��nk��KC�������<���x:�q�}G 0:�v�Q�$�j�B���� )��=7D���Y���rr̦˚,��h�:<^pP؄��v`6V�#�y)�r}�w�h�M��M�I $EI~���X�,��<t UP"װ4f1VRu��pJA�u�wy�V2�a�����}x�@�
�C�x�Q4�#�lS>�_�y�M���Y^�m2ҧg��$���=e���Ҁ�i������>�H$�-1�G�g�x�"��d2�\yۓX7�FgA�S�hFS[;?�۲��^��Tyv������������������Ʉmmlz����f_����[���+��a'k��w�@�E��=}�i��s5P��6L�8:2µL���B�cR]+`Rj��5�����D|�m��|ĹYF,%�`/�n���.N����j����#~�Ït����j����Q��P���2  @�.�����5����bv
	郍�;4�������¦t"}���|�0xX�8;'���Tk�>*�?�9^�˚���Wv!�,^���r�O^\)�·�pB����R���xyye�5TT>|������`x�T,�A[|��"~���+�:88 �&R��HPP��q��w+ ��PȯN�\�r�x�W�{������˭**-龫/8�wl��0�T���Nc������{��> �斖�YY�G(Mwwʘù�֬�����+<|��m^��	0?5� z 4(((F��0��2� ZW(!��AZݲI/_��  С�p����T�|�j4ONm-X��Җg�>�	~���Rmk�4�*k��b�W:E3<��1�l������<����o�Ù����˵��F:��@���������u0�ɤG�oO��N�'&&�E6�#D�R�������|"[��'�hьA�S�R�t�V�*�	.���謯ܤ^4���N[���؞iG���a�~(ƅ��s�n�����)Վ�낪��u��	������W���V���!�[>��L�������ܐ|��+!��ɩ)H�D��l�ܬ,�P2�1�wJ�_'��`1�j�	�x]n���N��&9�q���f.bv+�+���J{���5μ���S*��0�ȅ3��ӻƣ[5{o�9"9'8���WwY���B�%H�LSCC���<��3�+4>��Lօ �������1wr�A�:�Y��pk���?E��M��f�=����1HU�d9y�����n�S�߿�=�&f�U 8~YP�Ch#����H
}F�}�x�2֔��	D�6���|"�{)��o�����o�
���<���F0�еsx�5�3�w�xl���n!t��1�萸��CoŇ���څ���K|^5�
l��AQvvZ�N������'<gJ-iY=��;� ��yKO#���[�Y8���RfK����'þ���%]�w�mf��o�y����쑑�3'8�H��^���g7|�͙���4��(5�Q#�^���yy�G�:��d:��{�	�*E0�6��{�K0v�#sw�_�w��;/�d�z��`"��Ar�V�h$3m~�
SN��a�xG�-��uHIz�'s݂��2zO��^Hɇe6� ��3�c�{H8{~�Y�B��|D! �*gP�<F�5��{_j���8�@����"P2A6�bֹ�,��5�b�|iVś��[pB��Qr�'�27���7*��uT4{O
�D�x���ɕ��6�'�c��� ���g��qr��C+�(OH��mʎY���&4���%M>����d��j�WiE���K
�.S�7��PL���8��ۇ��[�gZ��n��1�����·wh��:��������L�P��o�3��� �ܫ����;�b�;�Mי���n����O3�������&��N�y�)���}��^l:Q�W��$Z+/D� ���ޤ 9�ΪO���}xi��ۺߢ�������h�x�}�RF�/��9>�[��?�4��C=�S�p���4�-��܆pX���n��/���DŦ�:Ăg���� zB�����TXJBHq�_@V�*Z��[Zyj�3E��vDw�Ŧ��G �z�r{j`�g��-��%�-���\W�w&���Ҁ�8���Cwg�#B�3�Y~�)�r��|f?�����O˴)�������{� ��P�T�Ҕ�m�ȡbO�X�z/R�b��c��{ͤ?�Z�h4����>���}}U`4�6W��j`�TU��;9>,=��� G/n��T���`�`�]Q�Ң�3�Z��4s����������������!����|�~�Ը�˂���{ISM-z�e����q{PH��ȌR�`����g����PN0�L(�~jo_1-��u�ζ��;~GC��#!Ε;7iJG2J��ˑN&�Saa�3�]�c�w������82��BK����Oթ����9���h��p���.�l[7�>���x�ծ��55Hq���+ �iH�5 yBK^�up���g���FZZ�P�"Y��E�'l5�j%a��c�����fݿ��Pڎ��"}'1$֢ݺE������72�����n�ś9�>�>�i8��B���
�e�"@	�hޮ�c�vT�k*���u��,߇�f��L�$�1�s�!�����=j�[�L^�7V�Q�J ����É|�Sk���g�����6:��(ࣷ�{�����g|�����\ /���K;��AK�zz�9#,�& ��.g��Чb^�$,թ�%e��I'�.��ׯq�0� )���s�K	dx]�U��폊)�D���R�;��h��^^��~��HG�F������V�X$ �ɏBUD7�A	F��R�	>@�x6}�����z���m�N\
|�ZWp"ɡ���I��E3)rH���W��g|����!� 9?�6������cc�%i��Hȳ���X��>�ՅG��]�����\Qy�z$W�Sr���#b�Y��V�L}��B����U�=$N�/K#�(I�n�mC����>$���k����Sy����ݫ
����--/�]2Ժ;� uK�������@|��zRq9MM5LJ�v�I�{oM��C�ZQY��VId��rv3�� �U�.G����qn����,n���C1���抉$���W�N�:hoA*��47OC7ůj֭�5�E�����'_�ЕRv��)�#X���-W��p�꺦l��[
��/%�`�ia#ԣQ{����Wu�e��J�p��MRR��!��'��V7m��CR3�G\����@X���[�>���O���SW`U��t�<�xX���tX�+,���MHD96�GŰ�[�� Ń'�L�����J�nd�D�ýX�H/\�
�~+�~[]�s�[���j�B~F�OD�逸��؊�ȓ?�lY�ᲃq成�=Qmy�/s�����55N:)w�B��yvW͌��z�vc�4Q�H��#iI'��5A�Z�W�6��{��L�.��U@�+'�ٛ���k�Fw��+�T�(@	b���9#T��f�/M�j{��*Z���������,=��ګI��P=���H�*���Z���f˓��^��_t�F��с�d��?�k~�h�<)ɋ�ia9,y�%S֮������n�m���u>��zӆ��R8Ru���1��3�)&d�~���Ց�[y���6�����{.3�je�V�}�|��@ ���k�B�5�r_��ӧ�HU���谸�S�7ɒ*����A��|M���k_:%"%�A~��6���ǈ��V��~[��N�&��Z��KIY.ˋ�k�'��Y�o���wp�@��ېB��x�8[_��q� �S���2���.�4����2w�p�f1��E�?KȪ��\ֲ�WS]��J��)WO�^oH��W����o'��V×��h�x ��lû�-{�{��}^��5�$�6�V����-|��q�(C�#gs"e����o�ΕΫ���s>���Eތ����%��d�G8<sg1����ߺs��b��e;C�����g�m~�j��ϬpR���4��<Djb�l�)6.n�~') ���]�-�G�����9�#XU�ü� �� %�����*��Z�\P�
���%�r�K����z@�v.h�`YYb�5�W�:sM���8[uL���"�#��B�V��}�!"�����?��������N���NM��a�Z�c�bM��]/��STbr�g-�2Q�:�{_m[��s+�s���+�4n"-uDq~�4�E�7��Tv�[[�ɼ�|)����1S�u�V�B�74��N�h���v���Y|`���q�u��[��"��᪓)��	S��0�{?��m��r��T#Z:�]��z�V%�����%^��}:�^��l�g�[ib\�D�֞Z���3���U!��.	6m�����Yݔ����ann^x��r�*����$��%���J�C�q,�E��FJ���BVn�S!�u��M(�FN8��o��[��9��؞H�#��O�w��Kr��٠�(���������R���((\	� ;5�R��3f!�JW^�ܸ�-�wj��-�g0+Gj�٪��ܠ<��`L�=�����A�D�%R3Ud��贺��)����@�3&�;��_��]>[�\?q�r�~�~�":Q��&J��A����t��=�q���jW){�zM�]���#:{��ʩ�!C�"��",�L%�w{{�f�k����l;@��F�����S9zH�h�uCBBx\�@\赨�����E[��\�9�[4�<x� ��{C�t!C����}��P;M�'֭�  3x���?;CtPf�ȟǓ^�(��7�w��W�|���w��t%�c��Q0��U��Ǵn���+�@�ͭ�/��;��}h�c&��v>��s!���4��M�s��	G)�e���iJ���ŵ�Z���1[C��F�K$g���.�1k�wx4��:h�`�=�m��ϳ���������U*c5��E8�4�w0�~�Q�L�a¸����� ?�b�t��a��j )��H��y3����
�-OʭƵ�,�EY�rɗ�
w�Z��5J�O�I�]�W4(m��ߺ=k��d8Fj�f����-*(Pn_�D'3=� K���4�I���u�\�����ESO���:@J�g�A�����:r�r��S��j�\�� 1�#�]Si�}���rߏӿe��K�y�t~����omu��^o���/��j��pPm�H��g����J�82�ͫ(̜�۫	[��)?5�l����%�Yk%g��j����ݴ|��{p";�O����f��8[gТ�0'G�]mE����qtf�t}�8����J��xxx��Uuu� �_��������ԧj��zL�|/2���}���>�&x5��sZ�W�B�g�}����O�EY=t�J6#���s�n���V�|�CF!�����Hq���.@*n�c�*��	ZliY7Y{�_H��|�x�ޔ�ib�eV��bI��N��M93#�4� �� _�1����mw�ɇ��._��#,|����m5!P�㘸�u�񜝝c�A�\Z\챐���K�11�tn�_�@��Q�!Y?o�����N�z����bS��6�[�ko��+��+���k�����Ma|�������R��O=�"��v��b��t�;�.,򮟚}�/1O��i�~zg$(���
Y�pG;XR�=����zT�}��Znn{SJ�=��q=PM9��!��'���	S�x�5c_�p�B|ݺ��
*���v=&������H�"yϨ��Fad!buX�{wb[��������@����?_0l��*����/Ūԉ9�?�ȋ�����H����o���Y*�*ٹ#���d��K��W�eo%t�{��$f�\���>��&+'l�<����ˬ�f`���q��/zc��G�cr��( �ⳟ.��Yg�-�&�ȩ��x5+Ñ����_i��)0���̾T'��%��'�[F���\�|��R�j�M���9��kcE����:����8�W/�����#�F��f�llj*=�Go.go��u#�q��qO=Pj��˻m~��r99��&�&�9=M���% "��vkE+N;o�|�=�ƴ��ѷ~s�uI���8�Ie��v. ���D�d��)�d��P������$�l��R���T��|�=��:���Z�^X�%���������{ID� W�����D���z����:����;Ϥ�v��zՊ�
�������n�Ր���������_pI��i����w(R0p+=]g����xJ��ԟ9�(�;g����Od#���{��d��W�H��t�=���"> �tʲ�_G=��r[myQ�]��[�����I��b>��N?q)~?������W�!��&���i}���7��p�w
cd�ǔ.U9���*X�B1�,�r�(�/{{PH�M���$m��*>d	�Pa�i���EU*�դԫI�S��:LW�,1����pÊY�0ӂ�o�o�D�6��>�S�@�GSsq�r��O� �͍'��H��W�͠^e��}&1�fP��ROdr�.�?��3�Ҁ:��Qq^�z��\q�S��r3o���25�c�wT�M$s����-�I�����M��v1��l��]�fKL.�֬K�e��O�A�d�����8�w` :������p�y4�������[��]�e�oO6�Y�҃fo�|�+��~�����/�2�r�(5TF[_|P��h��oб���� ��Qx�H1߃��N�>kk�DD�z/{7��Z[�K�+�m����� ��ׇ�6��"��p��
}ZyY��
)[�B�`�;���9�~���d���2��D8_�<Q=�bX��O�0��X�9��o?q} � z��!&�L��O�	U.@	�g��z�p	��,˙D���|7�n�'@��oD��x�x�ߝ�ŉ�ɯ�g�m��|�q�����g�����{;���U����8�jF	�"���1��U
�V���:Y'�pg�'�D�~U���=m~��}]�SȧUp��n�V�����¬��������۷H���]$�e�ꫝq���"L�=J��Jt�D��oD� �UL�{���h ܇�6��R�MW�5���o��y�*I;Y�Ք������N;���������mJp9>����`����<�
��3�v!�0n�n�1/��'��n�?̽wTT˶=�r�k��((�@R$K��Ar��AA���dԣ�( 9#H�"9�"Z�d����n~U��w����c����Uk�5�\k�]���x�A��F0?���B?��p�>%!���l�TE׈�l�^��w��*�!v��/�6��@q�x��}]xw-��Z��wD�X��^�#�$��CO]ͮx�H|⹚�_�_�N��G\�9K=�2�Cɦ�;s/�6��ͅ/�T��:�,ѷ�@K8&:w��yI�K�G��Sƣe	LS33e�F@(e����Xo�D��aUS�/����y�Ƈ��>ݍ�vA��?ٳ83??�� �Bl��+m�'��(v>�cYI'�>넫��:���������o` n���m�[/�T��v�\��:����Ļ}�W��d?��J!+����,Z�ru���͒��tW��N0D<̱,���M����������u2?�jxs��*������/��l3��O�b�e��(P��� J�jLM`��S%f�����:�P�^����ss+��iQ�� )�]���}2>z��9
6#y6�d����+��rkuOx���.6�\,ML����%#|�������
�����率cF�l�f���5��?��?�@���L�@.�X�@�y�ϕ�E��X�R����N�����Em��H�2ӹ�Wh�����E�N�P�����q������.{Q��1����̹'@��DK�����+��P�%���;]9���m��h����8�m��ҋ���n�i)-u�Y ��#t�G�<��e�)_֋�ݹψ��_����U���o��>��i^�ւ�m\��[���y�"�r�bq9�gMS���6�e_���kfq�,�ZMEW7��������)P6�e�����,�)SC��%�Ǔ�M��V*��P�;e7�[���!wsn:������ Ǘs�"g�/F�pk�GN����Ѱ��܎�:w���k����K'�*����pD��<��s2a�;�\�4�ǌ^�{W%'�΢]ԸjC��e5����6�4M���:4����^߄������O�|ic�RK��
�ԩ��\v^6���JkJ9�|yp%�X�3!;�p����M"���2P��I�	���j���7a��}EEG�����{�d}�#-2��0F�P-��סɮ����o�Ē�i���ܻ f8* ����l�TW�v�-g=����d�h7�Ժd�uG�����)Ij�/�1�^�>���j0,9o�ol�b�������%$��� {���T߀�.�=� G���A8�Q�%>�C��z�0����vVU����s�t��IU?�^��cf@a�I�bw�Yh<�l���,���#mˢ?v��7M&��w�R�.ix��J
nR��(������Y��*v!bJ����� �Žk�Ϋ(����ɮ���3Wڽ?�)��P��В�t��/\5���m� �M_��8E��u�1�
HZ�'{k�r��1Z6���:	Ӓ���9���H��$�p ����`��ͅ~�P�kxO�2�7p[�y�9m���FZMx�w? ��� ��fX�$M����则�%n=$�ifu��<@���Y�It������S'��' �̞,��u���"~���Q����M��@�uC��d��%Jȭ(F���@K��/ϰ��" �R��h2Y����=bt��i|>Q�?Rb_)\��q�HX�e}��V�9��=�<|W8jK�WJFO��=���wY���󻒽ڈՊԸۼ�_�� .��G��%�:
��BPb�1��=O�Qb>I��^_�$a�����B�*�%��5�P���� ;�\��-��m��l���L�g�m�yl�������|�`���j��w�J^NAa
����]Y�?.����\Jg�v_,�4R�Tz���eY4��p_��$�E+�~0ӕS͠9����лsYEL�91�`|n`��6h���a��w�a�+��Z�!c�a�5���ko-�.+�8�C%P9�Y-l��[]F��O�I^{���oE��=���=��#.����M�
6`�>~�����#J�N�_R�yY7n���;��2~���'K3��qN��*u������)G�4�^���_7��z���I��iX2�L��败�6󰓛z���P|�?��=��Ih�s�k�-�3I$�rt��ٹ3�!fbWt��+�@QX������W�
klL������4�����k$�.���T@����5�%�󿠷%��:��9y��O������Y��T������YRT�w�Ц&� A�������nf��Ѵ9*W���>|a`+ۙ���^�p�w������3�?�� �dV'�|Da�В�yN�4ũ��^���7�	�#h�33i�߾�
����o���_�˺/!��ٙ8�0?�,Mw���MN��{���7�B��f��p|���s�(��C���v�$]S��폯���J���+�h�}=�%c=7 �j�;r%�A�N-!+���p���uⱚuC�]s�!i�T���d��ﴪ�HR�×o?iK=Q:�DԖ&/o�D@����l��\�2]�X �'7(�ϱw�_?DOFi�&(>U�ϟ%�5ʗ�l��ګ�,@X<�Պ����j#�hy�w�O>�}8��C��V%���<�p!&fT��fc��-)��d|�� '"������tUDk�7k��G����E!�MP��N2HX]]]xC����P�~}:44�Ɋ��_9�2|�f��M���B.4��l�_�$,�72����Б����Z�Ί����8>{Y�u�
�������8K+����7\� � ,,V�;�y:���^gC���$����a�׾m����O /������Ve���_o��7���}����.���ٳ&������j��/nݺoUT�[DF�^�SQ]=�_@ �+E�[5��0 ��ֲ�3�]-B�Y�fX��@(l2��×�̯$�����_�̨07*��y�g���G�V�\����C����k�'){�>3�-@%-�f��W���7v���$���{��{�y#�51��a����� qS����|ޏ<��D�b@���%�g@Ut篻Tj��� ��KYk����Q55M?}�̤���4n��5���˵�/#h4�$�d3���v#���9e����̛�Y�~��v����j�+�� �͇��y,\�����Z��q�Vgg�6J�(֍�~���J��OJ��=�]��O���]�_�y�V�߶IXX�9Nvw��,�u5��?�d����)G ��[�����YwJ*��89���a������gώONL01���O���^�Z=���鱍����j}�ؾL^|��ӗ�i>�T�V�	&]	��_���%�̌8-#��P�0�{��&yy�����.{�ؗ���%W��b����v��Qa���gy�$tt��'jS����N�f:����.���?(������/����3δ� �g�u'p���� ��D|�y��_�����
h����R�W:l������E^3̋���#�s/�[�>��#���0�;��AeZc��R�֞��ӎ;��yP#lV����%UgX��Ek�t�H��y��iǙ!>C~��n���B�6${m�LF�,��R���]��j2w��,*3�6�S�GmZ�LI�yN�+���#�a��Q�@�r�x8��L�@���E����ٷ���a�pྖI%�p۔+�]`�cY�?7��ͯ��;�ę7"�iߘ"W��xO,�|t}�X�!��=��ä�@��k{D�mS�=�ϯVj��?���􃅦�i=K%�=�y_��	m���xVN��S�D=��k��oz`�Z{|T�l@@�٨�{��֩õ��Y�.UѝS����S*.�Ʊ
-������H;����O�j��_��U�.nx
3h�0�$�ŗ:�?��sw#������v�����5��6��EI7�� �1>K�����N��=>N�mf�JBs����6P���CC>����g�Z�s:���5��{�d����ș�S7����k�Hw�E��)L�������������
��㧆KSt���\���F���{��9=�"���}P� �V��~ġ��:�I+5�a�t���p�~�
Bܾ�)��5��a�Jfq�H�y����6.�&tͶ��Z�!L��~cᑪ��yw�d��A�o�(����z@��rI�CkI�J��& %'0nX�=	�;dx�*��wdj�/礇�VrS2j�?I�F�[�T�Q5�Q��}w�>�1��U�͹G�0�����JUQ�y��ǮX.��9;[֒��:�?�X᜿bk�E7���f��.�y�Z-��b�{/�<��S9]~�2����U����?{YԻg_�p�X]�֘���z�?�m�ֺ_`�^��s��SY 6�±��]�]v���qR��o< y�H�".����C`7�2xL=�0}G�Y����lN!�x��믤e�$�����!�^����������~7%����"�9���fJ�'e�bw����9]�ޣ�O,��]��Umc;����$u��L՟�+���ā�68޴��`�H��)>!ԡK�v�◦@0JSu{Q	�{���J�;�}�;�P�����ÙQᵊ�z�iXt��՝�ϝ��)o���0�>�!񘆆�������Z�z�h�<G/�uu�Bf�cL��>�,i�\K�ұ���'��6��ǖ�-�4�?���lZ�"^�\"��W�1p�A�y��T�,������W&`� �\Y�l��$	FjA Wa�U�p�3��L�|�}я��^�R�?+ş��i��7l��B�������d��4��mw<��{ש��s�ب����J�(�����f������v<�R֖�p����F�bt�v[�ZӴ�uWBG�f���@'.�n��y���N�|���?`���wс��ן����D[a�co�֑��|�������!w3*�O��Aչ�D;����[�3����#G�%fu���^��"�rA����ש�;ү�^��}���D^/MYvo�O�l�й�n��9if9��^�ſ�t��YP7�Qy|ڎ�VZ׎E6��㠻Jj�\j�`��J6Ze2���F
�x�N��-�	�·�>�\����Oa�eY|��B���N�]��J�Y��4�{C��h� ��d�A�e��v��O}՘�����A#O�D���w.s�o癚b�f^�/���9襀]�#�5g�@�H�h��d7��E}�/�DF�#}&Ks��񭭥+mE�w�Mؕ��`�O��rS����1�Ԥ{?���w˔Fl�%���#�i�e� ���Zl�����j�^'{��P2B <o
���@N�������É*��ᨈ�����J��Ph���[��"�Y�� �.ሥf��3¹��.����-rF)x.v���5���`e�?P���n�mdP�==�E��w �6�i��ʧl/���"#8LO�5��6�`E�7�0ۙ!d:�.��^�G#G���=Gq�~��e�
�X귳��R���ՊS�sf�4�,�iӍТ�΋Y�?������Urv:o�彍�l_xR�_l��}[Ͷ@h}[Co�8�̴<Re-ycd�����@�o��ܘ�m�l�M乁����R��)�6���ђ4����h�˶OTa��F9���8YD�H�����D�I����_��n�kn�ٴ�pu�W��xLV	}�Hƽr`����nRNH�ވݶ4�
��ָ���oF�'��L��:��{y��×�9��G�G�+X�'��FM ��x�8m�#T=C�6z�a�2^3�M��B�lXi:U_�#g�
���/�
��df���x�9N�LȂ��<yk�2-�˦b����e��G����M#L�ם�5�Ʀ^jl^�KF���F��ˬ�W�G�S���su7s�%^H��ձ�D�8�|��	��kؓK�XEl��]˚�G��+��	K����K������Zݴ��"Z�d��Ɛ���Ψ8���oF�X4z芭��ܐ��(9{Û�B�}��qw4l��&���4�5o���Η��V���9:��m�|*]$$~)�����s�N"��g��'����<q(���Л�BC�&��{�M����-���[Xې�G
"���)�^,�前 ����7k=�u]��oR^*ɋ쌽�,ΌQ��dc]��\,x���d�@�}W��|��;���Tr�=$�.�v����u�EW�c���AH�9�(,D��?ux��.`�>'��Ǭ����#��2���Q9�[0Z��R��I�?<��8"�cOhPO�6���~�'�s�ɉ��m����'|��Cb1h���'>7����:����?h��p�(���vhH&Y{C]ϟI���]���΀���lL8 �-h�&P�7�DG��5/yvh��Ж���r!@�f���2�mQî~l���M�8��ߌ!�	2�	*z�������|��l���/u�[�ts0vM�r ��"�&���@��ܼ4��d6_q�P��d�@��B.�F� N�D���ק���Q�ݍ�����; q>���V��k�(���1C�~aE�QQz��q�ۗq���۩Ω^49��sS�c��� 椠�j-�b��[o��ʴ�m��g�\���l�q�K,d�ta.ɷv��B�@z��i�B��>�]LD�W��cM a˻�h �"JW��z|q4�g�?uN��Q���T��*)c!M��s��X��>]�6�!���+��Q�5Bv$t��C�pn2�&.=���záMƃ9�W�k���M���_[�_ۼИc�?%e_CdYȀ���'g�>��y�<*��n�7S++����S9��T�%T�����dܕ�[Gp�&��C%��t��]�:�G�&!@��Cܪ �"�>t�d!W�dk�%_�ۃv=���0.2�a!ӠF���|#M0�<�Ĝt��$�K�n��2��|c�G[(�6�';�9�q�y5�,J�_�9�4y�`��!�&��A�3l��Vuz��:d�T���.c���͗�������+���'9�|Ӫ�����M{eeU�j>|8�4	��['�0���_����oƅ�V�&U����M��8��WcH��o�@��G����\ �7�n.��V
��|�NEF?FL^6��K��k�%	�H�(�
�;P��ܞ[0���e^D�)h����w����A�R�8����a��m�*���j��g}b�qϸi)A?گ����ţ_M0�������p�c髙�U:�����$lg���.MC��^D8���1�2Ѻ�I�f�]�UR�1[]YqG�I��u�%8��Y��Ռ��o͏�vƐ�1����tw0��
ht �_�����Ls<JV��u����ZM\�;B�a4�Rҁ!X7���T�<���I�����~� 7'U&T1�8��1�73��Sl��u�N�^�w%���kuUM��=v�K�yh�h�p��Ά��?��Mۄ����X:��n�6�[�156�ɕY�"|��Q88�U��$&il�rӷۢ�5��H*ሂ�F�Hnˑ��\�l����2��Tg�?3��K��ܚr*��LR��2G�*ߞntX(j�7�~�w��}\���X���-;Y������`��"c<tR�3�Wf��֢s�	V8��u��_��e��4��i@O`��&�]]:n�i���4W/z��\��</߸����R��(�߱�lx�T��j�aƢ	�~e�LȍO%���{u?u�I���]Ɩ�c������ߔ������ݜ��(C	'��uw��{��VÝ�q�ӞP��!=��oq�cP�zS�1�,9ǲ�\����f&���~ݞ	t�k9�FJ�0��b}�%�4#��:|�V���E1 UZ��>�k��MT�V��j�AR��g���i��|��P��5ť�z

,�WL���> 5�̗?�߬R�p�=��K:3}fxq ����Ú�.
&s���?�iS��6.�t�*J�=�p�������b�J0�ve���H N^�P�7�;
�K3��c
?��ȩ�2H������-���a�X��g��?w�͇���w��������(ݺ�;�l��53��r�����y����t�2�h�P�0_C���P8���L��*A6�/�f�F�T�Wo΀)u+1fp8NL\�V�G�9i) ����v\�v4�- ��W���0���(��d�*]"w����]Z�5���9��czR��-v�rwuj�C5S޼����1Y]v�rsz�d�����8(:�q���|��WJ1�7�:�T啿�[�{�o��44�,�� �#p�IFO�Q�E�dճ�r����<[��B��d�	�30$����d�X��zL�9n�;��N,��_wT�����=��ob��o>�Y��2_6�6�ڼm��BV܋ ��f��m�s�����'�pB��Z����3�@V'!�M�-ڝ@B�b�^����0��/@a/e-�:��X��M"���S�92U��*~dlQpd�{�:�0���ej���u�|�c	���A&B��FSUG�P9zl��a�`G^���@Y�
8�؃�!(�}r��3�&��I͍���zs5c6�ɦ3�������Z���g��Jq��P���y���2?�i���/C�k�+�K''�1G|U�FoLR@�s=MFE��9����Ӝ�q�)^6�@��.���C��-��3���-lq3���E"��<;���+F>��@���V\��Y��0����p��7�V�lj�qwz8��/��n�_��m�za���6 ��D�,17@���7��}|�k$�5��g'�o'(���YQV.�5y$,�l��bu�k�].�x�|Os�A�Q�K8����A��Ns�{�Kq ֦@P�t��4�d�����^�����r�Z��'�3�'ӏ�
<Q<��E1�i
W��E� ����3�����5�4����� ��� �
�g_�t(��3��f�m�����a�^��u����c�:�l�=��߽�k�x��w�pƓh�f����@��v撕:^2��q�!Ɛ��2��a!µ��yO"����W!)����'��s�Ut�����ț��g��0���;�|EA��Eoy��if��hq��3��tk�0�����1��u8�(wi�C -��<��c���A��Y z�0�#�cӍ3��>���t�L�F���?�:��U�Ze�,%\�Ԏ�͑.�H�~����f�??k>%���_��	��,���K��i�w���@��!e�Ќ{��J�_�������mRٰ��#���.
$��X����i�x����E�>�Ӿ��x�H�+����0����BR������
S�@�����'� O���+TQ��Ø8��T7�<&� YAmB���y�*�����������Ic�\ppc��r�'`�D=��Ӟ���y2���Ց��g48�����K�*�9ybA �+��b���/��!��<k�|�պ����&��%p�|϶�Y��w�j[6=O�\r^��]��#i
�+���O�ۡ���?Ì6b��d(S�i�..l���)���}4(��P`!31�H�c1��y�)\`DL�L�����LKUa�H��yC��3^��o�F������c�D7� `�����6�r6S��]n?8Q�P#��I;ľ$�/��:d�˗�UN+1�N����X�:Bg�v�����msV���O���m��v$�<a�>9�[����8�I� m���=��	DSV�]3P��9�uD�4�(�����Px4n���5��w~˯8KES���e�1��T��O�n�9�p����:RtS�@����w�i�w�7���Fv��� �u��|=N�ٿ�Ƀ�=j�E$)�7�8uw�&���e���q�)e�@,$��V�n��͓�!ǾM��G��t�F��\�pE���_���b��d9��uZ�0�>9��<�WX]�?�K�D{W��VW�v�Z�`����)�Nf�®��7�{��˜���{�3jp��5���`����z)I����T<�qf�
��w��|�mw�<Fk@�7, ��îl�O�6\8n%��d`Ny�j�� RT�P!�WR㻦�o����K8ȭ}�	��\�uS�_�����Gm���n&���T^K(`�l�c��_S������d6b��F�n�@F~R�50�vW��AB
ԍ���ۂq��ɷX�o���Ft�U�w"?�or�5��:��׷`~� �`��o��6��&I\�S�A�����0!����ݞ��0geh�pT��w@]qp�	��8�S�*�:��g����1�u����&�JH^<���_j	�ѣ\��_�	a���t_ ���"����n��L�ڊ�rB�� �É�3GB�%@3ϸ��8l�x�{��@�=��F��9�
9�b�����@�-�s5?�<J�c���!Q�f ��i�,�2�E��{k:Ku2扎2�m�/&OI�,u�2�n�!��
g��y�>n��π(�h��e��_0i���G!���uk��R���[����N�]�8T��緟�QA@"7��ư��'�{�\ެM3�X���B.]��%`��A�����Op'ջ��8{��\��h���Yao�t�aW����m��WYw����]	��%*���/\����f���`"��,�aY��,wnm�]:��g�ʷ��q1��΄AeF�o��|�:�pg>�t�[�3I����MX���ʓ�p�x��YS��kL��_�kPf�x�<3˜kKKe���y�8��:�P�n��|8X$=-8ʬL���*��A^����\�{�'p#�
��J%��Mse�v�����̰��I�Ɠ���F��ڪiH�Y������&���e�*�v�x�����l�D�q������/Y~xw�m����plv:sjz���$rx�����d�'�gLh�8pcǃ5���㔛}N.��q��q��a�fX|{�0���mt�a�H}�Ӵo�r�Y�r׎�����X�)]��8An4�D�����n�����⬫暟���Ȋ����W�4^�O\rLNV(9�#w��Lݾ$̣a�!��!��E����D�����Qh��4Ç�&�x�Vxsh��Y��e��/`Ws�"1��aNW�0 ̤0Ͷ���8�?	
�tq~9�VR11����r��>Y����m~-�I��<�z����_�k��{�k�Gpb\���'����c��?~LH�9 1'�55�IKTw7��F�z)��~�>������Ж�=�Ҿ���ny,Gf��[�(��n��_��� ��T�� ��&�+,�Y�,�c��j����r|3w��x>�j�������H��q ���Y�
��MA�7C���:::�Z9����޵WC p����`�[��i._(G�vG����7�wG�농�ĎJ��`����������l�2�*��zX,XXX\��GB�X˘Dv�EvE<�t�'���%;�b1��"��YFg$"N����ب��y���W���.yf��?������1O~��aֻ8yx���9HD�l���_�?sY�k��OlO�<Z��a�U[�>�SQCbbbҸ�Y�l��\�s��a۟��0�Gke��2��h�׏s����,s���@tΦD���z��z��E産�t���#.�E���� �,ݿ���p��X���W��,ⶐװJ�B�3�W6;;{|����m��C�~ZZZ�L�Rb��;l�滻���
�����o��X$+ݴv�\��މ��{����@�%赛�����}��j��ՀK�ǖ��Ѓ�q�9%�3o>g�U��L�Vϒ��mW��O��cH�6����ډ�u���.3	>w�j(^k���s���<����9����QV~Bbs`���#�}�i�����=$�Օ��ڹ#�� �v�~���v[s5hD�������x�l|���P�ӧO�۵B���������57?�'I�f(~�>\'H�cN����}$>ߢ����Nd9XT:E����5�c�:J�BW�<9�����م_SܹM��q�����FFI�/� ]�c�G�1��K�:����L����B��{bv�#ㄸ]�%t;� �P%㫳
^��a�p�m�2���s�Ή��^�vi��[���)T�epp$l>��r��+[��s�v���4+�1��V��1�M�iZ����pq����鮮.N��<�Ł��x�i��$���2>i������ ��q������f-�I��r�����M����Qt娌��~!4�}����Q���e�]��}����f�`be�H!遲���ߌ��S�m��_��.�ϑ��|�#;�K�l _��5�jY_e���E0,$Bx-��u��\q�=�Nl�?� x��B����l�������W�Y���I���JK�L�Go�n�VŴ�8��L�j#Fw�U]x�)I�ʭKG҄��u�t�^s�t�jhnRyy�����ɝ��U� ۟��L?#�h֑(�_bkHAI	�����:T]/23�,c��H�ɕ�B��V�'E�k����Xcz�'�����E�ۉ���=���4��E���9�����򠠠 �wT�uT����c��{'7�swvgN�:����Şb�K�9�;}ee�x��/_��k�F�a��8��e����s�CwX�a����������;��$���
��)�Άl��aέ�pt4n���:%z���|�U]N��w��גۨ��Qv\��2i1T�G�Vjw����r��yb�JɁ�^T��XM^ja!w4�����Z�G}>R80dt�&�ݭP���N����:�X@Spc��$^w����ӘGz��c���b�Gph�L��t��;�[$���>fN}-�ăik�ͺ��"P[w�W��d���`�F���i�i��V4�o��w��� TMMM�~�V,������3��X�rkR�vW�s'ܫt��/��Y�*�Tnh
	�q�TQ:�����P�3�מp�Q�$AC�[%�#bâ]4�9'bm|�
�UH�Whis��(y,��RN��3�Y�J'�طq���=������f^�dp��Dm�HjU�����#�$�@T|Z���y,�og"x�#�ӡwd��k��}����)�I�EN3@m����̜��Z�[�/)�J����q�,��Xa{��
������ҍ^���M�/ȧd�w��v�����x�������Nw�p�]� �f^��Ǻp[y�C�xl�p�OTtql��A�����b8S���K�z��K��|��#���i�����^�X$	��+���A�ߝ'Hм���W��{+�*���1�^<�\�(�Ъ���a^�͏_���=37	������Y��OB��嵫P�*����h�x
Ҽ<�d�^��^}V��ӷ�A8,22R�e�d���|d�j��aܵ�h~nnu%�Kp5�)?��@IQ�,>�`d��9��}�.��8�� �e	/�S6����ݳ7<h]-D���@^W��sqA���m�°T�r�m�855U�Ό|;7�!��ڦ�p;�ջ�pE?�ԋs@ڴ@v��,�e��i4Fܚ�^��Z�k��՘M"�R�hUnߣ��c���g|$獭���������|t�x�t	��t�*�M��]�5�����i����*~Gǔog��g�d�EM̱g�  �v�ݪ���ٌ�ʍhW{Bυ���GUl)���@���/|�'�ːe���:^�����o��c`b0�LCƦ��@�@����c��cB�5v\k�H\����$e��M-Q�J=��	=u�p��"k�"ʍ�G������4O�����5у�lJ�c�v�m�f܎�݁�m�#���uWt{� ��������s271���pb)))`b������R� ��M9��W&���������l8>�b� "�@��M��n�6�&�]Kb�`l�N�oۄ1�Ekȍ�^����C���"�Q��^��Ғ��i�X��n`�b/t��0o�R��?n&Ђ��Н�{�_@2�Jr#���ݷo��|�������ɵ_nɄ����g�Of=��S��˴X1�U�ck�C�Q1\�<e�_;���^�5F��>*?;/�$��Jl�]-[+.�Yj�������{���+TO_&xƈ�~i��0�b�YdMdz.3��F��q����} X~G�)�'Lt "�bW��E��ҟ�P�&wpp0���]���-��%�����hN ]N�A^Hv[�ܩ�z�P��h�%@�����OT��+�BE��2_�a���(Q*Q;��;a�I�`���v;O.�gR�kC�x#�2Q���K�~2*�5����^r�Z,���;p��D�8u���� �M��>O������z#̵���� ��T��.�%�����>�G�5\`G}�.��"���[��0d��3k�1������,�\C��r4V3++V�'����h����I,_�\�0�����Z�ͬ��_	�Fjt���SJ��O�=L�X����_V�]Y��%���EO�aǞ6Ԛ�ǣ�\*s�d,�����f)��-��×h�,@L�ХE/�#����8;��uP�$Q�-�Fq�lnZ��������W���RT����B�MC��6�**I�?��ZXV0K^"���<;Q�(y�fS�i�Z}�D*�ʠhyJ��?|���B�
������ ��E/!iH��N=����)��^R�T��,;�H9Ȝ�i�_C��{���J��f�����#���'����Tם��!ͤ�a��C1ϝ��;{=�7\�PX@��}w�~��z�xd��c���n���.�k|�sKH�V�%�p�@LM
|OZ��Q~	`��0m��լ�87V�|5���t"�;���G��R{Ǡ��oH��	��եu��l5�J�bn�M�1��2ۘ�w?�J��ݏ�>�0�Q�^�%�w��X���ݷ�0�?���1**J�43�
.lU�XӦSl�c���-�SAج�m4�}¨�f	a�HN����|��Fc* ��|�.A()+�XJg3����Ks��7UZ�m�.b��2?���:����XXX�;��q^9E�.v��ʣ
`���!Lllȝ+벧Qt�S����#w7����?�@]��z�'���B?��=�!��,!�	>Mש����齈�(c_<����
E��ýG�n^�_hXzCt�������̷�8q��1b�Dי�'����?X�[����a���=�m7V���N�C�rss��p��B';i�G�Z�Q�L���U��^_�cV �|ϸ]C��wj�v��G�H�!�7Vr�F�E�G��5��]����7�E(�{��� �Σӟ�n�� ��8����yN��W�V��������k��)�l*�ţ��eL��=d�4,������N6�D��\�ӈ���u ��ƭ�̈O�?��ၭ-��k��jzs�\�Ǻ���M��-���6��k� `�.0T��s:z���@IQO�&44�7~�7�1��V��j�m��K�z����oݻ�i��r{o@�d O���^V{��}(&L�{3�x����G���� �6�*A���i��
�19Q<�ZC^�p�(S�ۂ��n-������|��R�f<�!A+'p��^�o�:���[@��=-v�h��u�H��F�&U��T=�N̽����,��4�IwI�d�
�^426��2�.�Z6i;=7^咽DM�Z�T2�dk�px�'�@�'�YK��T�"��5�˝,׮�:������D��
��?ϰ4#uNk�N�Dο~%�W'�P_�f0~4������P�Q�v"ĥK����}����� ���ڵ������#qmƤB�A������r��^�y?mP��*XU5S��?�P[y0� ���t�IL��9o<o��M�%��HP}c
5,���2��x:v����%P4��1���˯�Q�^;k/���3¿Vп�I���73=]��m~!�D�&�΢Jo�_�	sΉ4/�?ox"��^⍯P�jj �b#9^�X�v�JW��_��xK�s�am�K_)ƗS��^�w�L����֯m���[*2mbV�����p0�'(�~d�W��\�$�uШ�1~.P�}��ff�߳�S L��@X�_C�5�<�W\F�)?��������D[o)y��|'u4������n�k�*��(���c�ySʢjq�q�9�yl��ĳ�mU����/���hc�Ƿ݇�`ܢ$��^`����1qG�kׅo�^�E�h��@>�d�z��ݨ}���J�j����wr�<�>�#QMYlݫ�f�_��vR��.+�6yE�u2�25��I-Z�5���y������'�����u_��%W�]�N�,<���C�3���s��|k'��O�A;��+;���������μ�2�Z|uƫ��+z���8�`�����3{=�� �I8�a�[�>^ڎ8O���M����2�`R/�����9�I�HY�n1�\*@���vuZ�L(�E$:�`�x%�W�GS~/v�͜ ^vm�h��ƍ:)��L�\��O�[_��
L�}p�Yi���C0���
��k�ɧ�D-z�u:]���L��O
.�,����>���������8��(m���k ��1=}hBK�ӎY7o��f!�.[i��)�A������rt)���}�|����h nc��Y>|�]#{�x]o_�n����~� ���v�-x&�D���gԸJ�oϩ4y�as����N���ɠr�L����e�/=͎�	�oDv���ّ��k?��܇�5]�=
k�l	�Q�XX��]+�+�F����yȁ;����Н'�>LT遏(�0��TJ8aH���9� JBC��Q?���b{��+[�-�š���d[^5�f�s�?����b��9�܁#]���!On���nwǻ��9l����,o�.�>}w0��_���Ł��n5�C��ybv����,��F7���=<�9��}�뺝H�A�N���`4Uuu�jO̅�j㶨Ɓq��1�e�� Z�`F�}�Ҿ?lU���~w����'=f>w��2��x2�D�����B��
�l�m���#/|�O�w*�'!Ѳ�zd�6��J����o&��-���@#s�
�C{�n'�@N��S���i-�L���ȵ�M��}
��׼���(ľ��,��0�{���0 "�UD�D��̳dH�NTm[y�� Һ}$@�C�KG
'����n���i�.R`��`_R�zXM����8��������"�b|q��ദ��4� s����F�ڨ���A�mN7v�E����K�&J��ag侴�ueF���O�	Td^?�����/���>\���q��>�p�h���.�'�9=�����Q�omĖDN�֘�s1�8��P�J}r�s�v�����I�������L�c�����u�W�.iXy�1�+��M�0�Z5����c9�R�54�<e~�β�;�Ґ%�	W~zg��7�(�.Um���^l@lQ�8��'�t����/>���r_�~��Dӻ֛�V�͸7�i:����ً�2�ʦ�5��z���;�[e��,�U<��l#Ǘ�&j�E���Vz�R�1�Z�E�ͺH�q�}�b��p���T��'Hh��R������1�L����/~2S-[�A����ݽ�Nse��Q���+�'�6�^'(���з	xu�����9ר����n����F�'��T�i)Ǹ�	)ȩJ��!�޶��ab]eǭk>�`ڕ"njj:��g� ٽ7����<O�(�z��j�������>��HO2��7M�s,���,�	�I�}@��!�SIW��p�.�
M�q&b�nFù������&���~w��5l���)��`�c�M�S�o|��ds�R��u�~��	g]\��p���x����gU����J}��������	)lT���Ue��8HH�ֹ�X�W�������������}�N�6J_h���5�Ƶ�[�N��� tz�պ���PUU��ifn>�(�#E�\�'{BԹ���yG�~̫c��%�����С�4�O����2���$K�j�U�b�:$j���;�c-z����4�`qp�l�ݘ���ǾbR�>\��6H::;wV�455u\g�W���&��)���:�₯�A�!�OF#r��-܈\9��Rɬ��?ʾ:*��^P�c�@@�[���F��.��N��N�.�����;���{���}�}k�Z��{���~���9'����[>��K��R�
�7�R�{ɚ��pW�=�7kV����pe�����O1a4��yD"x�xY�ևih�'��b���-�C��� �Z���)��+~<9������N��6�c���3�o(���..��8�<.�诏9���j��?��H2�SST1;_b@E������y4���v�U��M=�QV��!�F1����V�����t\���=I�����(.�r�4���]���xiw�螟�%W��gH�?�~�;��ˉ#l���bY��H��
fm�=���t�~�X-������x�+Im����|�}�A���I36�F�y�`��
�J�Vܝ?�Չ$���yH�Eu�Ҁ��|����Z
>ĥ�	����Ӆ�#3��^�X�K�D�,!���WFqo�}zi�8^f���{��!L�Aco{F#��6@���=����a�DFu��m�n�9��XT�R�k����dE��?�D��<�T��X�=~���� �&>�r��L ��JB ������l*�8���]��~��Dk"~g[���w��8Ƚ�E�:�l��5~��68�#���C 9��䫴4㔯I��w~x�S�y�zF`o~i,���	}���	����'2f����}�py��΢#0�|��9r�맃0�x�]����(�s��)T�������
T@�{T�k�G���=�⧮�	�1�L��~��F���bki���s�����;ӹ�;--������y�MU�&&�N��K>�/�ͼF��`��bP]z�),n��1˦3�PL��������X����v��g�$ɝ ���K�v�oo+LQ��>�6����D>;��Q�W5��O�����Q���.C<N�%uKf�YG��I9l�_P�ݻ���Pb2�ǵU���NwjoW僕���nr�+V�{r
�b����q,��c�aRo\�_i�}�=IR��}򾡥�ݘ����e�ͳ�p�zʩP��׽t
�N�C��b~?11��q�tņ�Av�����D��`������I�f	n��B���(����49�!�����[���mQ�]ulz[iAH��s����mx�rh��h��Iw�U�9�0{8s�됖�n���X$|>��р׻�i�����V���$�-�h-w����lt78�B�	��{߳�qG�,BED;:��s��.P���߬��G����D��ݵ�v�s.\�GMș/D��azq!����-�ta�k��"�2�t��q�*/gs����yo8�Ӂ�Ũ$M��}'A\0��A�U��[�gjͱ��������oÁ빧_V󢃼ff6'�����U�ƣ��K�h�J۶��`d;��@v�1��q!b�h����xY��d1��;�y�[ M*�������x��L�8�2�GR�䎳�cx,���(���h���/u�� Y���H�k?a^U�� ]8Z	��Z�H��v��3�ǭ�
,��6�+�	.��dt:[%i��\�l=is �_��8:�32��V'�XQ���ӤN�tq7���sK����ċ�ۉ#@^^\d�w��A�?:qվo�256�+��h<^�'��<� ���ZA@z߸��0�v�a���b�Ӡ�[c���H
.HD��7��c��GաҜSxP
���L�/o���ޕ�����q����>ɼGR�ᴴ��U���/ͺ�OU&i��oog�cIR������[]����� ��������/�y���P�8���Rd�[��uk�?eg���a���h� +ڍ�	vW������ގ�9��d�β��fh�ֹ�]y�a�J<V���A'̩N	� )5�v��ao��ս�*u)A/\��5~�-�0(\?}�j�ύ�����P!7KH���4 �r��tooo��o���;K�� e D���?��B,�kd?g�ڈ�ѽ��-�+����Se�ZtKw�<��/��������@�@�մ�J;@N�/�Q��S��h��MCAR�l�  �*���9]�l�\��LCI�*􊖖�_�~�9�hۤ����]�6PN�Q��A�%����IR���g��x2	���X��/I���d���A�
呪�ת�P��(��
Y��~�ID>d��x����I$+I.x��*-��� z�U\��B-<;�������x1<���A$�@�)IŲ>�;E[��7U��G��΋qg�ʇ�\�*�����/��:���n����۪�s�9��X`Tm=�3db;EZ����hMSX�4/:�h�F5�J�Q5#� �_����^^���"��3C��*�8�SR��A[�1�k�Ӎ.-���CU�,$<[Kz~�s��Pr��&��sV��;5.�z��JG�uwu�7l�Y�^�����\O(o����hD'�P�Hb8Vl'm�b�m�<}��Ư�;/�ʜ(�k<PH��6Z璻z���7JN���?
X�O#��{��~���.�~����\�����oGNm�s"�B��8��Hnt0�R�gV�6�-�vB�����-�̫�8..��E�X��p�`����Fn �w�ޞ�KPq� /���E�����}�ţǫ�{�A��z�K�ޢ������C���80���8^����7� �8b�N�+e>�ď@�f��XB�GEK%�����`����C��W��k�o�6?M/j�]�ԡO)O��hL���t�R�����x�P�w��l�P�	�?!h��'���y;�LMM,=N&�?�3-��7���.mD�W�N��3$��Ƌ�{���p���j�-^R\�<�EY�|�6YM���eGǷ�l8�����D/P�LD����a5�<	��>�M�U���L-�D�n^�Ի�ܼ���A����

�y��{�K`�H�8`�L�3|j�C��K"V:��Ǿz���Z"ל��h����6Y+-eVF9+�üb�b����}����B���Zi�.�HIK�ԗ���f@�숞���5��a�j\?Z��ɩ׀��0pXo�s���[A�R�m�D��?��ҁ�K��3��Ӑi�T���'X�PQm�O�NW���(���pX�uGP�	U�;�#yJV;��Ў ҡ� ����Gs3@zy�� ���o���v�M&"2�� ;=�](�	����B��9��A�V���Ư����68*W\<�[u]|�Z��n���l�>$"��7ع>N%�8�X?����{�S]��;��w�;i�a_�FY8���ZYI�U{��/�OlxvA���Y����E�.�>�Sæ��X����A��M"�a��o&V���7	p����!��}j(T��ߞZ��K5��:k͡�\~���7
-8Q�d%���& �P�r!���K��O�����#;Dl�6��M�#!TƐ
�/�K��3 ��h{�f��v莟wq��<�t/t�D���l�����1c+��e)t��4L�>xLr �n�t4����:�.aY�oG�7�\��<���o�_�nOO�߄.������d����-	C5`�a����4��j$jΦ{�g	��*0�;e�yI=�BTH�wf�����޵�s l��Q�
�׾(8K�σ�S�$y�t�ϭAx���d����a�'ՠ'Q~\}����ka��~%zЎ6?ܡ���#.�$��g �@|2RE���#p�lY>d���[Ծȶ	�1X�r��W�ջ ȨC�[$S���;�SSfn�*xP�Pd� �|»"l�NAϫ��O��+����Tb�dS^��<,����~�=�à��à�@�[ݻ��?#{X�FU�s+���>����o��/�vi8L�c�2� 4���U�9jcT��&�Í&'�@u]�!ujE;(p���FaU��8���X�6 �k��C7�b5/�-&!7�~S�"l�����\#��7k�B����I���5�0ĩ�d>#����3-�dL���1�S<|�r�V�ͳt,��b~f�FM{غ�Vp1!���`W���7��Bg���w���R����-��x{L��/���`���fš]�5�k%�&���ˠ/)qh\�}�� �VCҜ�)���X �4	ؕ�}�޺�X;��T����_�ᯉ�����H�M��e��P���Ο4i>�ᨺj�	���s-��̓zL2.fW|Ff��˶���8��|g��A`M�� S^q�FY/ݥ���^�Y	�>���L+��%O���w�	�4v۾xsF����َ��HZh��6����A9h��?����w�P+���3�z�"����ݵA 9Z �E��p&�Q���f���#�u�j9�!��+����A��ܫ��<���� ��q~

$ҁ7E�l��%��fCn���A�̰/ �L%Ǡ,)�)�4��i���MH ����9�V_�\�x�9���. %8ںpa?��R�2�n�2�&p������g  ��x��I�� ���"w"֏�O]�Z��U�< �uJI�VN#B�8v�����������d5X"QTV�w�Lp�@'i�)�[�>|��`>cuh����ŵ��#'7�o𓗃�� |5)O��Ld�d�2 �/�Qs8� P�@P�d�p��a`�g����j��>I��^��W�.l���KYi�V�p���ǧ����b��$IMyz}a^^ޘ���h�hQ9�~��71��i��~oޘ��x�	,�������
�^����1B%=�4��'s6F�b�\� �bl���� ���>z�0�2LϐP9�1�-�Hb��P`<�;���,�w�Kp3P$ƅZM_��+#��,�^�������`D�t9�N��N:���������{��%6��N�d�&���AsXjt[�rԌ�&A�n�C����r�U80��F+� �q��猫�W«�'��J���B��[ �{���@Lu��������"�	���b��t��	����T�d%E�6 ���O_V��>M��7| c c�O��
2w���}��@�����jO������T�~!�Fc�U���kEܘ-��@�	ďd5��q�� 0��� ��>1qI��N�	���4��@e��V��%���``c\�������#���'88%;�@�AK���#�n4���.���f�~�����\:�5��iL�ڕ���I�
�������-�������Z���A	�f��V�'啛����� ��3S�~Aq 7-���~ e0H���5���*V�6ߣ��2��t�L��$�A���Rf�ƹH�O�nG&oe+-��'wf�:����{�.��)Y~�b�݃��>'k��������5����QLZIeN�*��Ta ���^n$���ട������Ӄ��i�M�u�њ��3�@���X�٧� � \��\�9�m �p��yW:M� �G�V+keƒB��[��J�^k��s����bj�Q��py%���i���gacի��POE��̠������r6�n���6�n���i:-E1�`왿me�	@�����	�\�� �*�i��o��,bV�$�ܩ��~�k�p����aF��L#��@���E��@n����T���`#���ģ��,�Z;L�O`@0�Ouڷ:㧛���
X�fq�_�R�Lu����dHQ a%=-�i�M�l29��'a�]��$gZr��P2�VZZ������>.* ?:s�N C�/h��ZM��8�Ef7,�������z�(�Q&d�c:��I�x�j�(Ꞿ�w�
�mh�����1��C��7�/4O����R����.�&&�wM��e
\g}�%6�CT��`"fm�^C-�����ۊ�K)X�yo���A�8k�� �8�E�PHKo%�ؒ~���&�f��� 0��Ɠ-�"%��dff� ��IDʡ��zzz �Z��tһ0Ǚծ1��1���D��s�{��-d.I�8 ;�_	��w��\m�x<�79waV�Ţ�H�ck�k��0e*���4-� ��h��tHC���U�hύ1Ў��, �C���#h�5�����``���w!Ц:k�̑��(��޼�,`���2."�?�� ��,z�U��N�R�Q�<��د=?^�sv�6�e�uRR�U<9�Q��ičLO��h:���~������߆�Z�����"�}��KQ�����2���@Е�}�C�@cjb��##ZM���z����c��y=��T6%j�E�Π�b��������gq�%���������{Xb�6ȵ��>f\O��� �`�Ӯ����z>�4�W��"��ȱ������ı�=C�k�߱/�	�".�SKJXz��AV�\�Bg����e��ӫW�#|c��� ���b'�>N��c�D�'|���B����G�GV$��#�b&�	����+�Ʃ�K��C2777�����ܘ����_癞ӆ��#��	SFGG����D^N%h���ʅ�6���E5�q4��2�2& �hj5`j�q:�4�r�������������(({41K���M��k<CXRs4�~pAT��q��nC[�������ʅ��#�� �����+Eīz���9���w�3 �ϣB:���H@�H@�9`3Tޘ�;�6�ZL��Ow�%�܇ ��a����M����M=��7�����x4��D���2����J������B$©D޿�z��5�uq����_��e�c@���t���D�dL$�J�����cs��?�@@�f���E�g8e��| �Է�
�̮�Mޠa���Ke�|���X	ҋ��	������Lǒ����?~��L�l���`S�V�QL̘sJ�d���t�� ���$���y	]Z��� ����y�Y�[hӠ0�Y]�����6��y��_	&ڽo�^��y�_ɩ��KF)������<����+��JE����L4����c���<�F���{n]�iJ����;�ED�8�i��Ñ(A � �W.�=0��\����s�Ü�ZI���FD��g}��Z6�j���|�]!�q��&~5����SDX�c��\��~��b���8'�Z���J������7��A:�%�c��[�yJq�,��&�M�5�G�3 ��S�r=���9E4��
�l���C��8����j=i��s�o:���1L]���V;l�wgA.ic
�zy=e@]{��c�)s!�H�L��m��������μ�(����W���&��_��=��ޘ�!�ٮ�ɯ�H��S������{2�m^�Zɋ꥖H�OS����3ӬE�������	��{GdA�"�7Ƞ�F��F��?�f/�x���_~���;*-�X�|Ҫ7s�'�{��f����z�Fڷ�N��TС��][F��a��~��Y�`���]/{�`�A�?/��0�~LmaڵBW(���k�����UeX۸�N�c:��p���2�^.�ذy)p�pnu����v�WO����o�]8��x� �⨴}#� F_d����,^�b��g��q��l���P!u|�z�b�!��~͞�W�o�����l�,��'RS i�߼SX�O*�\�&Y�ޮp�t���q𒔔�O��(�%O�i�<�5֐�����h[�7��1@�y��((��-=a��bŦ��խ'.m,cM`8�'\�+�/bu�`j�ze�UW�]H1M��%���ȃ������U΅���"��'�1����#��6�ye}!)�^Z�������â��A���i�����p��X�W[J�OM���	��f��]D��yV�|�T�����(�!�镞�9k�T�ǴRri�џ6�Qp�����W	(fm: �K�1|�W�7yRn��.�K�8u�<L/3]:p�$Y�i��T�`0O���B�%ý�k`̣��t�[�1����~b\�����m�jU	�j���̔O�;��&`f
���ꁁ9�Z+.�ԟ!;4���?!8�#�@�A�(�}/�j�r������Ɯ�,d�=Q�@�?6v�6�*�&+\�.Y}����k�Zί����8'fL�1l9C�N앶m��L��Z�]V< ��v���.����oRT��	V�dVm8@�Z��0��hȧ�
�R���I�=݇Z��9�Loy�_���OFd���[K`6:|ۏd��^��cvb#�w�5�*&2z��_����
.�#�'�@	g�P�Ӱ�|���ڪ,�spL�G����u�����6%���j��<e���B	GN��VdZM��;%����'�޶�d"��ģ����\��LPKr��5P4]���=��w;��Y�]럏��@rWj͋�OS*���O5g��m�_v�+���'��eny�AA� �,N�`=��Q6e������r8HSꏒb�7�oWh5�s��z���1[��+������Qҥ���|��+�}lB�p��z�����(!\�˖D�[ה��f/�
T�z��f=#�Z��j�pq�,D4(��p5ڼ�t���|��L	|!n'8���r>?�����A5��F�6���ťK�b<�ItG��A�j�����Rp�&����S��ت28u:6��J�
�[���<�mL���*j9�@D�:��po��2 ^��3b��� ��L<��;ӛ��/����4�L��)�k��k���!y�*���%�ɑ����^z��
W�Tᵏ�!um���w�8�jkK�cL*Ρ��*t��C����ccw��K�G�#c��/�>K	&�g��Cv���j�?�-��N:������tmv��zh��i����f��\��~~�qj�ᙦ}E�܁�ɏIA�_�8|��(�X�qk��N�+�f�P�yY���i<r�.�����&�o<}]����G� _�������Z�0��D"�>҄%��-�
&˭2��2��UE�"I�v��*T�D�\�h@�ݙ�JSuK��:�y����"����'P��7�M�iɤc"*wp�9�@{�~�mf�c��3N�Ze6��𯯇��<�1*ac�c~J�Sux{��kNzMԹfa\Y�	����ڏ�Q>��_�B�Aʹ�����5"��t,#6oS�CS_>sJ�9R	����	�%�k��=!�M�о��N�޴�:�nrr��V:�E5�!��1��7v��k��H���d)&�o39ݞ3z-�&R�Ѩ&�S�TBH�>�����V���mI��䍈��{�3���b7�8�uϔ�����F�sCmE�������ő�-��L!��Qb���#R7��C��&5nx��v��Z�â��kr�a"�`ơ��OFm���B�h��k�_�&�6�����~��r;�m����W\?���0��xም��i��Ӓo��ɍ���IS��i!�*���PV~R�JܕE{��M�:�O�#r�t��3a(�l�C��w�Z�>,`���`�gs�w[�������\����=���L4T�l<��b�������w&����1��:��qf�ЙC�xgfz������GG��%s�=�Vp���]����ckWW�t���o�Ml�+���>��(��m����b�j-o�+"|�QhF���/D91�=�1��VO���5M�{���{YH3�&\	!�����`���q��\���9��8; ��^���p؞H��j�;Zv��n�����.��Aa{�1�q�SF�m����c�Z�Oڠ�]3���U��>��p�ٝ�ug�ȪF�[�!�= � 9��PX^2}�%����D"���tul�����B�owKn�(�-���6H���9P��P�M��Xu�`l��7��凮�6�`*��g=�V��*��ay�ݎ��YR]�`ƫc��{�4?!���7��IxB���!��WC�mP�7-��f󿧕���9�KI,��j�u�L�
~�v��n��:��d�u 	��+�h}�?y�qg�__G�FѾ�@Ӫ���2��l_���2s�VbŎő�������$���ݽ�����&�����=�Z�c�o3�ZH�?JG�/0�?Xxb=''2z�wnsk��]���@�it��,�η��RWo�\2n��vq2�"ԌY�	�x�4u��ac@�b���[֝�AN��|���zn0F�S�V��+G�Z	l���˅I��17�R���e�勳�tH�{E��#b��8Α�*�����B�U�|u�h+����w~���������mGN0U�~����.��ʔ�2�7`�CY�$DD��ɵ�����n��G{ү��$��>3�N^�e'}/����p���wo�7��7�·^�-N �p%SAWڭ��俖�)�trσiyhЩ������{���k� ��>s%����?"0��Ƃ������G�i{�gv̇}�59����6tm��)ũ��:�m�pw�'_-�Xߕ9AF�]���5�מ�N���|}t�]�F��u2�}��*����<��0n'J@�ȉ��5gJWe�~ܨ	jH�<2®�����/�:�i7���x��m;�p}�	�U��E��|�ؒ󀑢Ì[�V�c�R��*��
u����2�~b��*�m�qQ��Q߉̚�l�`l���&�2���+�?-�1�/,�"���.Zo8���4?	=�����&�K�J<(ެ�xH��-�G�nc&:���Zؚ��Y��99���e���]�ځ=Cv0�� �Z#�"��m�mx�4���K0~��8i�S��>[*aO�JmH�;�}]5�ӌ�E�nHL��0��<�F�W]�9��z����!2⏱���s��JXH*�ۇ<	��Is6Woj��-�q�8��R�R�Ȗ���21q��#ǖ�����c˻����XXV��ٮ�����;��XN��$�͚;�-��U��X�Ol�-��<�2��3m�Fa.i-�3��^h�xO��K����z�/~����35gǖ!v�fqJs#��4��^�<r�Oj���o��
�ƍ�&Z�~X4�+�N�u���z@���K���N<9���\�?"k�38d%Mv��U���T�bg.��m��W������9âmE"e[lƢ�):�IX,;�g����d�Y-uy��V+WV��W6n{��8��:U+,,�E��W�m(wߙM���x����{RpR쳪p�p�Wr^6�lH\1�g�fƲ	9i��0��g|�fłԕ�g��?�r�U����@lǂ(��W˓�b�{[���C�1��W��Xj�D��Y���d36�Z��ڪ�3�Q�\�3s0D~n$3�v�>�QQ����怊,r�*=��q��]i�$%��k�)}6+�B'�#�PV<>��|��-ru�Yr�7�b�����n5�F-ֈ>���*�����V��F��m�GT���>����~���� �w��#r�r�k���^<g?N�D9�ؙ� G)����C\0��ؖ6���ki��fbFk�M*���D��8=}���Bn����՝V�H}6�P���,jרD����h�~���gu-�LE��%������08ߙ�Ht�k��M��=���HyIٱ� ��RHrH�[ t� �k����;���4խd�U��Aҟ,ז���b��G|�z�n/oߎ)xFJ-�r"B�O�3fe�:-vp|;Nd �8CIDk�k�k/2\�vb%��n00֘�+6D<�$�9��%�b���Dn�7��8T3��Σ�9��x������+���QO�O
�,�]xT;��+�a�]����ϵ���tC���!��8B$�����2#��o���,��lI]��0���Nn�dpj�F�R��(�O���ď�{���)>]���S۰�J���f_��,-���T����3���[�G	�� 7�^���v~��X�"4�,k�������`��@eT���M�#'.<?���k��N�oZ ���G.��1�b� ��j�c5�L
�v�o�Ww4�1W�#�5<���Yk�8������,��d�E������V�]�#g�e_Ѫ~�rti:�*�aT~Z�:Ms�|��`cb�`�h���}�������Ǉ$�O��B��S��uV-^�M~[ؠc�'����3[�l���;��	ɋ�vad���u?�-kb��S�jq�~[T����� ���4�p8-Y㖐��;���.@�ɲ��RT�t�\���/���4,�@�����]���D�%Q�^X�S�|w�E�����)�����EJD������^��}��|�!��Isz3G�W'����
�V�^T	�+��J߄��{bb!���y�3�@�$����������c�`���A�x��!���8��Ǩ�ݲV�&0��3Sɛ��&ngJK�Ԁw,��8�V�?����*F�X�����-ڗ>��U%t������9�k
M��n��Ԣ���c�L�D�ˢz���ɷ�|\��6\�� �Ӵ�zMǵ��7
y������GJR]�hu"����#o��!ڮ"���Jr�`K�K�"v��[��>��2޻���]�z���"�kL4�}�L���=�?I6�$�d%���
O~\�*@�"jc}������*6`4�c�����T��nV�

z��L �l���=�1�]�oHw����ɴ�e^z�s�A�����O�Ղ��P����+?c�E����.�Τ�����xS{��+�d1�����VU���s����0N��ه��j I��|�:T�ῑ�]+^l�����A�Rc���pt1�I�2�
T�|�wG��ihl�T�`���%e	����߿���Z:Y�?׎��uo7��d4���(�#�Vw��U��J�ER���0|�'�� �D�Eܼ�*��#�:in%|�tz���}r��
,���Z\"�w���v|���i�9=�{Sx�:�`8���{��99iZ=��b�^�L�x�p�&�����O&m�^�p�2�S'���D�[��,]� r��{�Y�XՔ]]�@�0�_�h��L�q��x�!���)�K��h�zݙ��
�������g s�Tnx�X��ײE0��|����/������������݊�V����P�HHe0Cy��x�	!�yٜu/c�r���%��ok��v�������r��ߵ��;*�o�6��U�5y�J�xR5q4���훨����Q�f�p��4����u�0�G �5k�7�(��EC]��)K)�d_�n�kB�y�ɤW�����Q?!���E��шOg����D�\���ŷ2��t��h{��80;Ns;�%�uޟ�}@t���R1�a�˨��r�t�̨[�bw������ok��Ω��U��1�t%��������:|*�BgC����O��n�<���v�<�I
����i� �1Wj [	5�a���O4�*|c��~�b�~~�ls���~�E��k�?rTK�l�3c����h���Z �U"$�8�lh�0j#K���т�}�B�a_Ử�#�1�ʽ�t&]��c�=��f��@A�&ڳ�۠�kG�m�B\ă�7�]�Tζ-�V�t!��O��t��f��`#��j��t��׽���(	���	z%�w!�3�����*86�Zit��f#q�ڕ�`�ė�y*3�����c������E����L���e��ʠC6���n��g�Ќ�l�������*ԝ�u=ph춬�u-�<MX�E��%�@�:h]7��F�f5[�s����ʢZ���o:|���z�%w���n446x���p��$*Sa08��To��k��4� �N�34��墪s�g�Oq]nt��,\4�����޳�C~;/O�T9߶(,�f���̤.�?�̠����Ĭm0%$e���42������;����\	�1&����I�D�	���*�Q�ho֜��{�D�$�N~p۞��_}�ϟ�r�q�W���uLME[�4�W6y�n�nt������� .���FOoE@�}/�EϬD��XҕD�O��\���]���uѝ��* �������B�ۛ6��>l���^���߁ ��C���a��Ʈ��*`)'�n��(��zOOC:W��ȵ�@	s��#}R?B�����jphJ�[��ivDN)M�0;lsg#���TR���sI�Ñ��k�miut)~W���чs~���	�4<˼������������[=P����A��I���ŏ�x��Dr�( 8�^%�,�{�TS��*�f:�${\�&�G��pI�ǕA�^Rz�Ŗq'ͤ\S��Z1A�j�ϩչ7�4^&�د�6q��l#��
�����U��G�[�t���5vr%���X�ǽi� a�y)ۃ�-�����??�v�����k��r�tw����?۴QB�H<����p(��,�]��ۮ��xrQq���1Ǔ��d���".�r1��^O� ��C�|v�IQ�q��&�Rc�'����^b3��?
��c�N&ȫ���¤�8�h Ⱥ���nC+~�A��Y{�ͳ���GvtnZ��5O�<��3�U��u�N�+= �� �*l��{.�e�l~��o�_��1�
	�]�1wv>P��Q7�x���� �Ѳ��(��!�S�f���.b������aċ�v���G�q����G�Y�� B��V�������6�'l��B.���}y�f�<)3�(6�Y'�����7!�U0k�F�v����Zd_	�����>�*b�y�����#i(�<Z�kY}�v$�!�;��CS��z��P��2��4}y��C����
�ے��,F20��Շ�^�<޷��)OH���'�������=kd�#Q1�}<J֬�>']��V��
7��xò�v+�,?�,9��?9G����)��)ү����s�,t"ˣ�5��T��w���iڵ�M�&��b2p�/���1?�A�/�����������l ]q�_|��*��N�C@��A�Sp8C�)�6�nx���oʆ�\���V�,|G��s_�(�j9d�`�_��=���n⇝��D@��k�D�s�d��i�����ݶs<^�Gϐ��|1S��t)�O�Oǅ��0w#�׸�s��Qd���v������A����c�?{����EThN�chm��3h���_��\E�Ҋ���7bցN~��������Y����(�8Q>�`͉QK�@�hw�����	�ӝ�O�M�OQ����i#����"�r����,������_�L�e����L�FaVAf��ʛ���0�&�]���f�G�v6�c�jզ����	ў� ��{�T�g�����Y�Ky!_B������z�z��w����`�ǝ��ć����
͜����,J�'��ǳ38.6}-3)vWd�Y��Yb�6��Vd�!Z����Op�9l��������m��/��o&�_��S��#���]���d�w��+���� mܟ�r��ȼv�����RUN�6ۈ��8�'�
|1�i���߯ �><��&���(���6��N�9'E<� ���_[y����~E�+�$]��vC^��h�]��S��c�Nm��b��⦊���.
�L쎔�i_p.�O�G!d}�VG����'O76
�r�ǆ�#.�֒��ZİfWOlq���Y�@v�0d{�y�O@,����h%Se��;����bM�l#���n[���ζ�!7�ۥ�P�u{mp��4,��lI���.�K�u%OB������J�!e��kM��z�]���+7����&Q��y����B�璂|������ﶬ@V��4̷1�ܰ�K��IU��b<��C���
�k���=6+�o�j��<B88����F���Unt�9��G��Z���ћD����/kd˸D�n�Ҕ���x`�,/v]�e�;�A�A ;�pV���������l�Q���V�Z����}���p6�̪��G�i(���?+XtI#���Q��`h�8܉r���yL���/m�����y�5)n������a�����UeQ�z���[L��m)����7BΦ�ˍõ�;��kp��!yZm3G�)���Z�^�g<3K?�%̓db����n9	�2��L���1a����c%Sd���J�4eƅ�n1�ȥ�1	'�0�~O���������r��=0n��� $-7�ſ�9����|R#Q�['�0�ʔ_[��!K�x��r�,P���]C��ɭF�[3[&�w�I�N��ii�*I�F&����<�y��'�3 CO�s�]5���3��ZIa}��69+�1bq�OB�5�'V��/��(B�yu���s��mO9��n~}ދ�����󙙊��3x;���_[��1����M1��:[k�H����̯�lU����>K�e�ˊ�F����A��<.�ض}�H^p�W��v�X�H�3+=	���f��k�tC�;Aɔ����V�g��E<��V�˒#�j�3Z֢��x�RةQ�k�Q��S���W�=m��\�j���~=W̓zf���p鬭'e���O�~�O{�73`�s�;>1��1�*g��/7��b��^��M�<yN	�/<�����祺�?�B�~h�g��Q%�����Ns�o�o�Q�(�~�!���/ːR�[:	'�=�`�(�r8Ӱ�:�(��I�͜]�C�QF�I�UM-Ua�M>���OJ]i���u*���I�Tp�d=	t�(Ő����G�$u �D��G���|���QX}�x�_�+��!��y����\!�0®(w�0�#.�-2qg��'�����%E�Li[3�>��t$� ��|~'ՄR����;�QlK^�u[:��5�ѭ�����P��GjZɓ�f�";}v�|�m�Pgt����)x�Cq;��w%�,��8��Gw%�q��8�zh�w����o��[u��1����e���ˁG�T�Ϧ6�G����"�]�y*M���y$��`l"wl��bϽ�t�J����L���d8�ia�!#3���=�'�?w��Mv����'z6=ƒɋ^�B%IH�8o�n�8)T��e
0)�E�C!`�^^UN(�?u#Ȍ5�
�_�rD	D���oJ����#���F�
�e_��4��3j峸������&��Djx�=#��p� pB�,��	f�_!����QXef.z3(C	��eD$�˴@֊ �,ZN��~�	6a�zh����������I>  ĕ������*40��Vi����?���f3�9�+KAG���ߣ>�Q}�6��~C}v<�J���U�����w,��������[�+J�H�/��o�Y[���kd_Y�/~��-�|���~dx=���U��W1c#n{�%
K$jE��9h�t<2Y'�WP��{�ﯡ����#A�)m��Eݲ-�-p��)a�X���f��|��	�/e�[�߁G�rt��Һ���E��y�{J��}~U[rw��hc��x�7~.����?��M�V��=��pM�����0e���l'T�<CH'h������u7F�<�W<�x��a��dҽ�㨫����*����T�IgED�J	J�AB��WE�.]:H�n�B�Dj� B%� ߹xyޟ�����br�̙s��:s��1}�4q�����C,1_.'���M<c�D2���Oπ��<�hae�)u����v ��IzL������F�4�)���_t��ȕD�}[�k�6�B!�T��&��/��;lQ�v�뗽�t�h�sS�ɯB�'���O\��7��&���������j�s6-A�Uo���u�7]Ώ�[a_�sq�:��d�8������Tu��W�&'��uՃ�Y�����m:�tr��w�:^�j���B��J}w$|���/O�c�����4t��� A���Fg�æGݻ��/���A�Y�B:���	?��Wsh�,���|�O����`���H���sv�ɨ$�$L����Zn�N�����H4�z�,WN�z �)�Yd��vEA؏gUg��ˍ-H��x7��tfp��$��_;qz�^�)��wS�[�rT��V�W	8"G�!��WF�w�(�@~�}�	�)����ʳ���Z ?O_�t�a'���e����*��1�c�-���.���r��}q2N|�}y~�(��Wq�Ni��Z����$#"�߼�0x�ks�i��F�0���^�T��]
*&\J�����he} �qif���K냫�d��f�.�.}�+�*k4ig�d*�l������ �VW�����M��k�E`7�l���h���S�	m'z~QTGN����]n�:���1r��@�@;���$�����_&ku�/���;�Π�ѽ���+�t�$oַ�����iD���c	�y��[�}x\	����瀃;+������K�����tWf?4��-�ҽ�YK��3�jc�x�s4�yo:��}�=�[W����E��l ��j`�:��W�a(:p���Rnя<��iW�*M6yi���MmE�;�n@�\� �H�q��\8K��S�C8l��U۷�Ǡ�z��ӉP��h�l���5��^�Y(r��F����Te]����K�0�Y?)m���^��率���9�i�ژ��뒮c�F������
^��sR�[iXOWX�Q0�b�/ϼ�p��G�l�?�Y\b������ �X����_�&��m�%H�����>+��}�jn�~V�~��F�3���(���D�C3��lu��$2խMER0AJ^+�ё�8o��U1t �`ݮa��:�穽�v�N�i�|e��閘���~�� �>�Ǌ���>�TK�T�����օ�t���s,Wi�.�ʯ�$�q0��o�����\W�n���1�?i�b����fg�Eq�!�����`��Ս�+\�::-δ�q���O��#k���v;�]t0�k�?������(l�0�O^����m��.�n���2864/�r�����TO�WM��Ik�w(���ۍ��[Zy�._���f��¡4�J��-��&�	��Y��������}��-a��{��,�T�`�ʶ�I?{��C�o�٫BNv_V���;A�}=l�%:w�`y3ñ��ŃJ��:���`g7���&���]gu����
v�>�+���F�j�<L�=�N�笛�lI��W�Rc�Е܃A�Zm��5B��v0��G��j� 8sY�x;t�%�������d��N@��.[���,0Q� �*�/�!��~���4��q��6úI��g�K��P�V���j/h���s=���^E�'���Z�GGc��gǬ)�/�F x|��_��馫�O��Ё�Og�o^�|�H�)+������2[1��D�i�;�0��J�*z���'���a,��	�{���0�m	c�[W���ͳ/𕚤�ؤ,-��cb8Ulg�Zk=}�%��,�N�n�����f	��Jo���\�ġ�@���0#�o}��/	^6��O
 r̚��V܂����#$�����ט�`�K�Jǎו^\��Y�rB��C�D��r�c��'���m�"�8�O�U�=��~ �#z���僸�o��@���8�;��d��&�^Ԋ�����=�᫝ʰ��G��v2k�[�9�� y����i�FBģf���(�����z}]��;r�X1阂ם�i�׀�!�*㈲���|�q�4"y�, l�����*����]LX�\~���m���N���_\����r@��p�}����`�HMǣ��M�J�*b�_��=F�+�%�Ux}��B��A �>JfGػ6ALJ�V��~��Ά�t��7TgGt͏�,�s�1)*]�\6��쫙 ̭���t��#�������A]Q4�8�W�Z[[u�k��ir��F�.�ww�$�;��a��e���l��w*�4�O��Rޕ���0-lQU��*?#�p����&��s�/5�^b��z�*3�K��w����
��T`�[��nV/ܧ�A� v�h��&��nv�U��Ȼ:�Up,`����k��
�Ba_]h=*�)���.~݀d��M�.�&|���Uu�\�����l���PX�����脌\���o��O�H��X\�Y���H<NCII	��y�^��5 8̚�����C�a7 ���u7�!���!7�zt���7�>�nf �y�+W#�3��rƭ�W/f's������'�åk�����uwC�p�~������)� 1���h�H�:�`�� �n�I"2�2~3������.#��I�����F�}�uٝ�q0�e����^<������g�3�4]��楤܄�v=~�a����d:L�c���$�R�%�;]G�p(!#�˥�pd31f�}�V��sY'�������L|X�j�z���ex��	�5-��&552}�m�tө@¼��6,�2q�M��b�~@�i�P�-;~�ڿx4�_F �M�������ć'��2,��f��=����O��[�׿�>x-CT7�������i2z�_8�z	�}%bB2Ew�7�y���/�B�����t@O���_�~7����/�k2�d=��=�dG�1�(@V6��T�f�B*an#��z9�/ߥ���K�v���l�G�\�"1��U�5*8.�3��r]��'��K:�W��Ƥ�>����S
�X4l�h�1�����1A;�g�\��<��7���߭ߍ����*�8��mᓓ���0y�\��*��ۛ�T+>(��(��Dy���,��o�%���/�U��]�p�x���L�G �x[������3"|�)"O�_�+�K{���8{�-�!)�"nk�����f*� h�f����@b��!mrL�srs�ʇ2���^��0�叽fݢ�4�)u��e���g"R�-f�~٫��/�X͔�|t��.�@��+j�#çt���l��wbw���l��]�56��2%��Zy��6��m+X�!�.8ő	 � ����T"3�U ����v�h���,D������3QQv���n`�{�v�Z�0�%�t���R���W9V.�V+x�Sz��h�nrҰhgsuvu2nX$�K[�c9,��左�Ʊ��u�ܟ�VR.�H���S���-f�'�.��-r!er�l��	���y��0��;��0���Μ��I�!7�̔�z�D�A77F�i
ރ�'��	�3��N���2�i�8�� �*Rw�������u���?���v��;�9�,��n<���3�#��}����M��������j5�����A9��=��C镕2j=&(����e�'O�퍔kv�P�[�w�JF�ok�yH^P*�땭�U˽��l�Y��V�TA���FJ�� �^���r�l��T��lݮnm�_Z�h��=��I=҄[F�� `��w}��t�J+@2#�~ -41�--
�X�U�T��=Y�Lqv6�ߧ�Ta��5B\�ș�����2���wGW�p�b����k6g�����]���q(B�Z@@@Tn��t�{ڠ�������]VTƴ^�7*��+6Rnkl/Hn����©]i�~Tn�=zר\���-�Q����+��Anm��!F:Z%��a��u�u]�y��jS��s���ع���>t7~��YZh�"��~�����ׂy�PƺI��(��|����S��Km^ړO-LML��X~!䀽�����cG^x�x~�I����b�6w}q��P�k��k��Ǐp�����|�W����p�P���A^ݼ�`����L�u�?�;������j�l_�җIN�oO�$|c����I4�8��SUHr�'��l�$��y��v�v��5�K+*��ߋ�PG��,�cW��_x��~�-�2¢�b([Օ�5�F�̸���W�a��sǋ�h����>hr,�U��=BO��oW`���S��<]���#��5�㘤��_��t�l =��,��}��GMb��^�_B�*(��j=�����jW`��l�;	]:t�s�V;&�J�Z@��}'�|E�T:������6��BH�|�h��H���s?cOz�i��1��N��!��R,? u�j@�w��uQ.�������yZ�Nۀٌ6�CF	����wc�nI�jvC�RK-�ε��w��Μ��9�̗�o���L5���|��<�4S��Wu�5�`e��
��VIl	������nܙ��cٴ����L�]��R F}�40�Rs���O�B~}1'ے*j���ZJ�=["W�Y����q�6n����v@u���s�����X ��ia�6�a��sNsC�}s��}������"l��=�	ٚ}���/�N�M�*���WӅ|��U�!��O^V��fp�&esR�������F�2����=,wLȯ���<�8mAI��H��B��V���w;0Dyg����D�ƣb����B�mo�pr&v�����q��
 zSb�A�5ͫ;<���z�5ވ�6�=x�?���[i����;v��Ы�S��(nA�o��: 7���I@�Mm��\����,����U���SG�Y)-�m[C��`��D���K�~0�4��^U�?���5����ra嚻�Q-�
�4��U*�����7��wxr䵝�+e���%1y�!�V\O����Q;��>v�baS}%ı,M`��c�ce��n|���o�K�fI��9+��|.�c��v�����M+G���d�Q���1����QMt���Px
���o��ǏM�q����	�����*/�R�J�M�x��@6�۰�%��Gq���3�'�YVM;5��LM��s��{.%�◫���m����7��ݎG;|��?����2v��������/ΛGZH>���K�3#ڪ��~lJjJ,��o�������M�p1�Ƿg��3��C�	N�Ya�jjj�%/�.��~l��b�7�����^iM����w������i�Q8=�� Μ0$^`��Z(��X��CIJH̛��ӓ�q���Č�dQ�)Uق������5�=��-i���KL T;�ʜR�;���>�V���1'i-?��9ױ���-�]�����f[48]�m��JI�KRF&a^k;@�«���3<%����Ro�����t�X\�{��i�A>1�O��>Й<�1�Lm�w{ǭ��-tAb\3ڄ�0��:�~��b�GI�j�d���+Ű��":���r$�&g�&���3����}_���c_�<������2�C^4Rhd��0Z�rH�YYΩW�d�6l�v�����k�}���V����[�W���݌d=wn*9lll�K����C�@7�,��PG �g����PKtu�ʞV�Yl!7MdD
(u"ѳ�I�M���YgX���H�L��I2������R����A�i����$�D�����O����=<u���rw��b��r�ތ�z�2b*	�	{	,p�|�WGKYU�����nŭ4�<Gk��j^�W��ѷ=,K�Okj�9�>!�7.Q�CZ��,&fI�)>5;�w��B&JT&g "�����8#m�ӥ90��߷z�����vR?�?��l�d��K̳H\2Z�j�튖p?��9�\�9�;#P�NK����D
b�(�v(t���O�GVo�^V1W\���l@Pv^�c*O�Y{H�����U��H��#+����&�v��?��{z"rz0�g�08_K�ʻ^ĳ�� u��z{���ߠ�$�
�Y[�Y��5T�*�}��5g:��1���{�т�ETy��m��X�$O,�آ%
*B������z��+�{=X�޸�5�@�#�]��9����1M֪��᠛}GϤf�_n���nOʳ|��Iq�-��Fջ��k��<�J�7q�
)�2_t^k�Q�u�L>��Qs7��c\N�0,;���궢�#!���#(I�p[o��Y()��Y����@�Ы.�x��{T�;�F�8��W��旡���H�J�b	�5�����V����沁)6�2W������Ħ]�e5R�K�����^�n	KHH zBtM|�%���פF��T�Y���E���%�B�0�����n�27b
�����D�!0I�h�O�[u,�ٻi��"��xc�ccxPni��t�Y:o���f��Uo��5�缵>��g?͡�\�8`�>Ojx1���>H�a6�[�e4��g�P3�0��JC�T&̆������n�qv���j[`�g�y6�|r�P�tn�v���c�o���F��mmm�-������<1�EV�D�q֑���D薾0�.6��w�	���9ۭ�`��;�nM���qF?=�g>��h�j�1�Y����yEb;��l�n�xתeE?�LtB�a�2�o�����<Gq)S��b�y�6�Ƹ�ZO�b�Ȩ_�ـ��SeQ�dM������kݏM��t�Y��L%Qk��M�?�8~B����x���M��}�._�������k=(��tmAtW�<������^�[��CԔm��ޞd�����p8�A~gɇ�Hj1���Xzmv���~9�<� ������*F�d�96�8&�ב�TΝ4J/�*/�7�>�E�V�U���m�Pߙ �U�TT��H��dG�F�m؂�h���짼��Uvf�^{[_��t��Z�7_-���O��������
�:����P�l%�J�����0�ø9]���dsP�p:p��� B[��sI�k��Q��ND�.����|\v�S<�p��� � �$3BC�aa�"O�dUеh��:Q�J��˞9�-��,�$B9��`c�a0z�;MU���j�jr�+��of��z/T�g���������'��j�8�2ǡX��������\��H��|%^v�)�����M��՟iF��f��C,���Ӥ�xd%W����D�(&9��_��qt��Y���#�n��R1��){v���g��g�%��<�;�ځ���%�[���LO�F�u����}�� ��I}L>�K��9�Y�0}&�>ǂ�p;��|��:;xHu[����e@9���{�,D0���
܈l*i��m��i�HGI���r8�6 �X�c���h%iQ�"U=q|&1z�ˑ*a�2�#��k#IP����*$Ȗ;+�K�pn�����X��$��T4��� W�����|@���H�=�"y 'ǥۅDs�>E�D��f�f� ��2����OU,d��* �	}4!9;^rh˾�v�0K��sń�2�)A����\�qn�:�dYru�n�����c����C�Y�'''�P1�<�����*Ae��^��:��^���IJ&	�M���w$\�&�%T�Z��^��K#V��oN�p��,�޾b��+�Br���5����1re���F.a�Rp��ׯ�'���}����.�c-�4ຘ�j�IbWӳjt[�J�0�;��T1Z�<���i�c�3���B#��%��g��6���b�61�D�]~Sk�����2T�c�<�������d��=��"4��Wi��R	؞X�<a�~�)l2�r�r���̝����»(�JR/���t�N&��3aD>t�`���}�*M�*L'���,4�"�y	~T�%Ҁ4��g��N���U��ER[[r��Ź�"��xi�F'H#ևܭ�k�}H���%�'�'�j}�L�G����.������Ġچ���\�o��b3x�X6z� Qߑ+if�~���sR���%:�[�+���M�g�JmZ��������3����h���pg��j�v~�r��'D�32�%���gڪ}��hI�����At�n�֤��eu�������f��sZ�:|Q�4�@��:{xH$3U�~�_�O&�15�����՜m���WϏ��;�����;��K��;�s�A����^�7��7����&T%
�j�7�6�%J�"e���l4�>W�\ (��a�!����nL?�U��/L%������e>��>Q&�{� �����j��lLgn\��E��*W�{6!�����Q]���\�P<;�F��ʫ���-����		�r�)�w�z������v޷���egr���928���Bvt�7�,l�����N��Α H�� 㪮����c(:�'�y�"L�xΐ��p��YU0�rdy>QhCE��c0��^t"���sۑ��)�tT�L�m�+qf�j�_f�G���v��_���u�z�D��I~H>�2����?Ҩ5`�N/����8�&����"g�;K��.!�kM�T�4Gls��u����B�l��T��lu5\���_��:m�d�"_S���>�qM�cKs�Q��۱�X|����J3��8�^Y����L��l$Q�`��؛?�R./;��������+r�y0~� �3�:Z�MK���e�>?|�p T�4��;U�WI���n��n'IH
U�����o���@ê�]NL?B�~�(Jd��s��_H�#�|=�B�%�v�Uk���?	'^Ř/�+����c�}�5���S��˟7dy�Xz�[���L<��1��GZ�>�%
�O����xK���/�;��2��{yRӲ�3��2�X�����x^nN"Ԭ3\�yˉ>��Xb�7%0��D��M��6���]i��V"z5T^znZ���^��k�I�┌�#�)�n��/p��m�>ݝ�6>$��iQ�~/�'��)�;��&�ؚ�qi���������Q��lZ��em���(�7����(��B=��zz윤����~	�r���n)����!m�1 �������$�wRs��R
��Z��J"W�&�g��� =���*KX񃒉�Dm�U�o�y�R�3����m5�zv����޳�4�4�U$}�=Z!��!T���N�$�7r��B,�Sv&J�J��́��ܩ~�uԽɉ��3���Lq9џ8|g0�9�3��9�_Bp��!��h�(�_��.�U�<� H�r#�̞0����Pl�Xt	�
��#� �Z(H������ezO۹@ �E�������/�=�F�w����d����=�3訛������,vR��i�~ߙ��CN1+J�oO �뻤]nX���@�n�q�AZ%PY����A�-:�v�{ڊ�x{�C�M!L��.i�
Kž6fä�
�o&�i�Ƨ��s�Y�`�p�\~�1�Y��iV�2��M�����!�"����hUM[��q���%�͇<�Q�.i�v��1]Q��!7*�����=�m���e��~Nq�����!cyL��*�e��p�DT���}�v�Dz�u4��Z�J��m�K�J�L>o/�	�V� ��1D[�t4��f�ϥ㻾ejm�+~��뗏B
�O��a�+J�<1[�i{��\d�揦����@�:�5܄ML������~@H�k� qpF�(
��i6t�w{7����C�M�1)��C�1�ZA�ҥ���i$Y	�e$����` ��3λ������F~v�E hb��B�8W&*8����ɛ|v�T��](99rR�n\zZf��*�2-������ĖIX]]��.x'9K5i0�i�2��DJ�D.m*��/Q0de���¯���`}��}v]X�Ў��'��Ǣ���͈�p��H�h�>]ZZ���Vjx��[�]�S��iI;q�hgυ"��O�~��_�
Z�z|��S��[�UhC���8OI9VD̸I�����_�]V*
D��Q �]<�p�����I����7P�o�#.Ck�@|� ����֖�9J�� �
.G���n��3��q��m�ȋ]�Qk�d�A5����~_�S;�h�_�'G�y�J�)���N�?��Bn&�K�}`�be)U�Bư�@�V&���[f�ʌ�p1��C�ǁ3%^s����PN�{��*�Xxi�j'��!�.��b7{��G��*ہf<�v4��`P����D��7���sϳǾf��v?��M�.K$:��5��,jbFn(J)�BR�J�&O<!ї۸�3t-�-dpQ� �ek!�`hf"j8=Չ�aQ׳�f��9����o�&�y��Y���&r7X���K6�ި�L6�;@���&	������eq �4��+�d(������=�j��9�u�%�r�}z쳆`K;���?�unv�k��t�s�kS�fu%jm	$�_�7��9��վ��JBpr[��.%�g@4�z���x���s��]���n�]������r���tc�12m��Y�M���74��툪7rq�A�慨@�)�mЂ@�k�� %
x%�����$�=l�R�-5��аˑ�Exࢷ'��^�	H1�5�rXڲhWwB�erҍX�a���nk���G�v[�(�"ۂ�fP��7��*�1R�~��1H��	�/��p�jB��� .�\o�z7��>&����GW�;��h���y�Ѿ��=Gk�����P/3s\����2 ��5�T�`'}����{�@��1~jƾ��0�*4?}��Q�u�\"d&X��;��{�C�N��,��a����4b��d��u���A�h �ZR��x�ڧ�<3LX0�L�`�{�D��� ��E~*M�G�4<�
ĵ) =6�T��ȹL]���z����v>��K���'�#��'�n���>��]ZU�K�Z�v��������ِ*�_�[1�t!�J� �W�r"�<�� �BYi�c
���� ��_Ly$�A�\���n�l���e�Ӫn���5Y0N�Ά�y��D;�Zk�C��`��p�Qe����	%e�0ݜ&�7��}>��վtJ_�mޜ5Zm�8�[s�����R�k��]����a��d�A���`�r[���W�\�P���k�K>6,.����h9KX������A���AG��lm��`��e%&�+�N�����M�_��k��= �	>���/��R�ݵkoM^;q�j�R�%� �A>�)��ùL}ِ�u`�Ì`zW�.�6LuxcP�O~�i��!����~gO�2�J_����_���}K=1�\FL�l��5q�p�bd�o����>;�n�~!��{�OM+����%@�^-Uh���OOl��VݏJm� � �)2�Fz��r�i��Z��@�2K��hW�#�I��׈(q&63�gg@��Ci8T�t�]_��"8ug l�"�W�	xD�f:Ż���3}����~���b鳪�$���8�f"�2N��	����g���þ�ЍA�P��]��i _- _���Y<��$ew�YŝWo���L���TG�ϖucD���d���1Q3�v�B��C��[�ò']��=K���2�r��0�ɐ��SjyL䄆(wWnGL��1u�� 1r�9�I%��3l�	{@)����A�ԎQ�/5��J�0��Y��#�!��p�Q���Hj���P��%i��#��v�y�v[��2dX�����1�S�%�T��7��ӏ�" [�nH���ڥ���^�pt,c�c�_,�`��Z�0�߳}y��`�;1w��������`K� �@�c��]9$J����7�`F���Wn�~m�"kl-���©�#hnY��#/�4�Ux�%��]S(���c -Or쬊��j��fE$��w�wŗY���A�&+>�,Rf�E�K�!���P�]�ҳ/xM�>'�F^�{�~�k��9uOɞ>�d]I4I؎o��x��9�V��ܮ�hS?|wd@�j�̶�k G}qB�8�Uj���L�q���#u�v�{\����C�˓�4P���ż����B�c����ӛ�x]h~.�`���J��2ွ��9$7�L�IL5��G��\�o���P��gj������z����l�c323�o�>����Jʒ\����˃��,��u��^�XN�W�K����?����h]S���x�Db(-K�ޡ�]<�=6�
�R�;52�ӚPB5�x��M�v�F�=�	�[I5(|��~o4��ȝ�Y�ԏ��.Yj��ww$��Y�?�>Z��Abqdgȑ+7o�z�r�ʩ�S�e�䆏Ys� �M�K&��ʇ唦Ծ�Lhn!ќ�y����~�5$	��a�Զ�x&//�e����ߗ�w�=e�K�f� ��S��1AMh�fPs`����f��~u�����,�>/ e`�U��5��S�3Fa\��wgg/���]���Dul�{~�X?�Ez�w�^����[E0�V����y8� �&X��DJ4�_1KF�ti==J� M{�յg�"�R^�V U���$lE��6�L
�>c~���H85=h1��[�'��*�v���t���n�z��)1 ) `R-��ٕ��^����Ԑ��Jנ��:hu}�_^�f1�BI91�m�x�0 CO���>U��^(��3lԽ��=����{ȄNCeee��l-�Ђ�;�b6X��J�O;[O��h�ĭ�<X^.S�'����&���E6p��ԑ.#�3&�s	��Op�g>-���~��a�("�;���9��Ώ/M��i{{o�����a;��ڑ�F��_���x�N�Ўd�e��U:��8�E�)��8������%����9���>D��L�є�&'>�ݰ�8�M�X���?��)���>��*.f���E�j�!�BU�۟��B�s1yh8��ں� ��i�y�~SR~z���lR�`���ZLڝ�/�����#- ���1���c�N�-�&nL��dк����\�>R5�g9<����Nd�]�:���	R���rMu�H�4,�s������q2^��#I�i�~�}�gM0�#������+��+����$ƍ���줌���$���$l$���i!@���#�� = 6��Q:r������^I��l�{��r�G���J�Ԥ5����[|�q���m�2���	���B�a�%�ZX(Q��٦�ZPe)��E�!��r3_�i9%U�Zj6�/)od3���`pw���X�^pl�	��]��Y�5#�6�E����S<w��w��I[��[�V���S72
�����ho�=�� ϗ3�:�>�\s��b󦰔T~�_Ϡ5$�"8�+�X�~���|�E�?����������~2^���3z��N�6�Ա��O��u��)����}Z�P�>��la�p��Z�m�_�֟b�e�h���i/���+���=�ӥ �ձb:#�,���j�{zM�<�������}��x.����������N�6����rˡ�Ko᭵�
�OlS���NF�Ğ�[���g'����w�����[VWW����T�P�ؼ�|���2C��93��b����j�)��//���_�K:_NMM�qtDC���\��_<����<�Vbr��X���1��y9�/9E�-.:%�u6���Pմ%b���ǖ�W�dWu���9M����*o1�U��x��2�fFʩ���5F�Ц�A��e�8!�;RiʯE��{�D� p>���Ǐ�~�r�$R���	�i��`���xt���ϗ1&o�~-t��z��I4�}6D~ǃ�¿��!�Q�2��3gơf�"�n_������x��:��%�� ͈s�j�&���Y�?/�'Y�S�b(���+p�o��bdG��J���]��,r�(>"��W�[|<Ж$��Bq�c�'�r��o�����6R�<)�V���DT����P�[z�`1�$~2���	,ԸE�W8MX��ʊ�@ٮ�<;D,��]#�`�������vh�yx��ٹ�i�{����}�:ٜ��!�C�6�
.��������x�w���#��j���!�nZ_��YS�{}_��Q0Ǧ�r��sz5�ݤr���u�}mv5�5,'�Wrsrr���������oZ&�d������]?ʺ�|���+!�T,���:��{i�s��暍:�=X�`)�Ơq����|�N%5Q��=[�3��[��1L� �);�V���_�
VI��[Db�-o��5hK�nN�ᄁ�������J�?��.l�&_�c���V�c|���^n��W+��S��|z�S�����O�Є?c�����7qD������y��ښ�c��K������A쟘c�Ρ	8e�lu�W'�*���P��B��FȢI���#��g�D���sFf ���l�v|�9O��6���W�!�����Ib���9&۶����-͏ݶ;��K|yy9vn��3�rC��{526>�׿�"F�RCz&����D�{�*�;y2�u���$˓�/���IzW���P6i��9�}WR$+�{�YZ	W�XZa��M��ua�w��ӱ�/~-t��kmU_#�~�ɨ��D��������:a?2�f���\�k��wM�ϐ�l�;%���6!���4T$XLRo_aE<�G�"ot�/_�E�Z�aº A9������2Qr?�������L����+�w�ݨ��_l��L��ƯV�Eb��}=8�x�=\����Ɩ�����? R��{��PNX|n��z_�	ԶV�t���3���}C�b8t�ѭ'�Sy��4�CD�o?��#���-�Ժ*�u��ω������=�^yJfF�X/g��s����3������@9\~Z'�����l�s�(;���g�r����n`u��]�=Z��gBR�v��">��;�ŋTA���l��9!v�0���������7����:㊀��+�@�J,C���o��e�c@Q#��������
���CX�tss{�Ƹ/t�@7��L��4�Ғ	moo
���6���
1����Dg��eA�_A�����M2��Aj�������j��&��}���`����6�&���)t�ٙ��N]�W��_u�x�S���N��ǹ�Mb��_���=5�.�����'롽� ��ȉ0(�����q���=�mT��l��`f�J�����������7�7��M-Sk)�a��O��&���L��(ݳc�I�܂G�����t��7(}�΍�3E�Q��V'�C��Vg��?�x�����߳�`>m`�������|�՝xƄ;��w����.�*��/}s:1�&�J[��C'���U&�-�|j����$���-4��.�&1j��$T��"~�Z���� h���ׯ��d��A�0��������à��\g��.`��J����x��s�j�c��v4swr���ޛ�:t���5�#Ф=������ç/�@�����m;-����ĝ���k��'55�������-����5�;_g�?�K����x�l��E�MGG��򣽯�
=A�D�|kLY�UR+���+���P|�W��v����m���,�@����s/r����KK�ߌ'�BB^���W��-$��Y��K�|���:��g��mq�/����;a�J�c0��7U 7bqm>i�z��V��m���Ǯw����Y����A%ї�0~��k��7W�L�X�����O��9wmVY~�tO�^jﶣ ����/���DT��� ��D��Ɍ��#��D��Ћ��u�Y:34Zl�A�r���M�IЇ5u�;ߡ\����C�l�������Dog���_/#PәI��,O�\�u'$�Ͳצ����\�4\b|��'3�.l�m����w8�]pCT	N��:��KKK�L�G�~��&bkg�&�3�*٦`��O���,|_e�5'g5W�E�z�U��v�%�x]��}P�K�_��.���@��zz&Eµ������dÉ���6��Z�^r��%op�6R(��|lx�LF�0��� ~�DO˹j2A��}_T�!�6S�1~@�/E21��zK.h�G���Q�|�c��@M �m�Y%�}��db��������3)�?�31�0!5�]�l�����?��ά�HWCD=�����x�����w��U��Id#]]�	~E�xori"\k��P_�+���`6ր� Iכֿ%I�,`f%++�|� /��{��	�,�)��\^^^�>CF����Yl�`�>��u5G�Y٪i���T��Y���+l`���'h6@����9���]���R��Ĺg����M��K_�C��?;=�Z�l��SK^{-��zŷ��Z8�bVʌ�~-�E�K�@\k����V##�y6������eα��Xz�$i�����h�]J9|�k5Z���=�}N�}��J���b�I���O�س�9�s�عf��3U����;5�kB'�6F���G|��A�6����-%&���A�8Yq��3�m�����X�ǻ{J�(��o1>�"�q����*�	��F�0�	d�����=~ iA�������n��l^QH{�T_6�����m����� �:߀l
����=ON^��4�<8������g��&�HRϙ�!��0�#/D��zoL}x���0�����`�����o�>�z��{�	�@g�]`�A5V`@����|f iu=�l
�R�
w]�������fw�@q^K��;e����ډʴ禪�N�8*�!�c8r��`�%��o,Z�pR������YqQ�Q���8�[�%��Z�3X�w�����2�����|m��%j���	m"S���o�� ��O��h)>&ÈY������к��f�/�:��F>�8
2����ӯ���,~1R��r�[�i�z�ީ�����RGs
�?�>�砼-��mA��:�/���Lp3�7��1��Cj1	�^���k� e�:66�����:�
�s�#~��`8��ܬ	�ZzA��������ռ��#~��Ǎ����	�>�9[ gyo��|�]�OS	wf{vq��օILR�,��ٽ*�z�T0^����>�c�~F�(|��އ(��	cu��\B����g ��r��l�^�v�)�\���б:#�-�դɍ~lux��<�&ծ��2+?��
LPI������o����+-{/�]���3p�Ԑ�Sb6>RFd��D�]Me��/Іn�����b{__�,��zVxP��j��c�ɞt<2�J�����u1V��r7�mbO���y�;�{�u(�j�w� Ғ�A���!P�	:?�E�F{���?����9(v������,o��Ю��dA�S1���o������rR�&Ɂo|4���c��Ӽ��Ҩ6vV+�k�H���
Y�.���"s��8	���@�[�B�g�
���{ �C��x�,�F�݋g��wQ=_����ZK)��D.���Q��� �@���)/��:h�@x��]ڮ��Af��-�^��؋�m��4��c�f>����.���l�!_���c�����F�������
L����l���W'u�2#���3^����Ϸ��_�5<�X�m���5v��w�3���".�Q�͡�I#����Ng��`/Pv�p&�����+�a�Q�sy/}N�i��������1R~��S�6���J~/r�VF�3Pô9
l�/K��8���j�b/R*��Z����BK���S�lu�v����]T7�2(-�{�0��J��g�9�ˑ.�A�������H��Zp��J�p)l��GL@�e�>��P�{���u4�8��B�ޛKX<l�'�u�������{�yAMT�ݺz��M���۳)E��#;�Y�x�u�z;���x���T�O3�zG���o���z2WP^��C�	��=�q���>�։��ڒ%�'��t��68 �u��e��rj��ݾה�
�Tʣ�6@���w����dojY������"�+����D����|�.u˫	K!�l�=�8�=�*9�����dT�9���Ç���l��AOG��m�W���i4�)i��S�W"�T�]M���������۬y�V��.��(�S]"��[(��8��޻���B��2��$I��BZ�Z+���JTō�����fi�T��I8��H���?I���P��Ɠ���c�-��Z��a�(�@DB�CZi�nPRZrhT��n�$��A%F�`e�a�n��������%�x�l�X�^������31BJ$���ƽ��Hg��������I[�7%�掸�`�_8��Ғ�#�� �r��4�	�b;�~x8(7)����Z��V�O��:�_s��!11W�>�Uu��l�c��t��;��*ãS<�Ӛ���5�'4��^�ϾS���'�f}��R
ibg��s���	vR�����L� 	�[!;��J��I
�Vήf��I�S_�ǝ�D�vUf���	��h�����j��u������h��6h���e���D��r�F[�C���5nv����J�%���)�p�(�2�8"��/M[?>�"Sd*q?_b{�,T�ض������ez�(H�>?��Y6��]�����r���O8?�� ���Kxjr�bǓ'߂�an�U����,����gv�4���q�~[R��R��q�����9wt n�܏�q����Z�6�֒��y�>�~ڸ����R�;+�{ �F�x�P�J�>2ho:[�2���f��ô�:��2c�E�F*	83�l{3��M���ن1&�u�7�WQ��E	Ѻ19� �v�׈F��%���'�[D��sz�ģN' |�ǛZt8:c��c�v���`�N?�;ڽvҢj�S����E�=���g= u�Je�8�Ѡ�&�Q�-�E��&�ə�o�{��;��QY�����������W��X��=׈#�X�L#F��L���0E:��������.���M�4���']ϩ��.or0<������(�!�c�-�m?���C�nh�{�6p	�y�?��Ъt��g������4�ӇL��O���ޙm����^,��zt�joNu[U�a1$��{+�uz�	)5�N{��(����M�<�ڐ���{�ȇLy� q��z��׿����UD�X�{L�"��JA��v%7�G��]��gk*�DM�Q��="%d
~���s��9�ۘ�e�п�����f`���O =$%##S��61�v�}�Ȇ�� � ����KQ�eq1bfo���v�}�~��4?[GvEF�~��`~n2B�9���`�8Uؓ�7�uDb��z�i ��	�KU_7-����\U����Y�|�y ڋdfa�ilBrqW9-t�6����qm]ݢХYc�L�}ι8R��@�`����a������|> 	*}�t����;.Bs;���c`t�ifؼq)�fv���(
���}bbuky�L,��)u��b�Pr9�Z��[��rN��iWTD^�A&ehhX�cf�4���̼�3���6�Z;vȸ<�N��Z���w���j���yh����V�O��P�r��)�)λ�)ej�^��Y{��$��S�z٭4�J�O���Ylqvm�m��� % 1Z�>���aIU!���U��8�L&����->�f�(�����ZV~�z���hl�]����n%��V�<p]Hl��W��o4xeh��P��{Tફn"���P�� ��g�g�j�K��-���3:�Z'P���[:�6y���T�2���[�D"����Y��e��T�yWtu1>��TB�H�Z3��x�"O��� Gy�:aZR�?8�
�ѫ��7��y ��Y!&��������>GGJ��陑E��	c�6��}	Q��C{��=ʢ A�@QeUK��t���9^�2A%O:����`��FL����/�	Z�h�͝�یfES'���rt ��G9��Xc��) .&�ieo_ ����n�b�'��9�~����sw8,~����O����@N�tG����x���Լ��\�cߓ��i����r�����e�|�h���5�&����?�F���<�Ydu�-bS�ڬR�yU�E�η�!��PY��^F���}s�~1�op:U���f-�c��Q�!�qYa/����(eb��_u0O��L_D}1��T2�ݑV@�-�MDI<�0d~���M�"?�Y
@��X�eȠb��C��a�H���I��;�>�bAL��d	_U�����k^�4h��ǁ��n���f~$��{�I��7լ8�ޚ�z�:����P�~E�=���[J�~�vb6P��dԘ���Ϙ̵�r:7���}`�흾F�(�_��8A�cp�QU�����[������U��-�j���!��0��m��$��<q�`���Y }��cP��sw���:y����1�i��nM60�'�+pA���@X��e5&^���[���(B��ZG�yQ��'�x�rRטXe������i�ǯ�r����ȁ�4w�g=��p=j��a8JC~d�kk�b���"���&��pj�%�r����;��1?֓��z�t�A�ᾊ�L]o:L&����K�1��22���"K�x$���� ��Xf����d�	����>.�|���39K�%>+W�&�����sG�9��]����b(Z��C�]�F��(R�C/�U_�W�wˤ�I�3}n�l��t~f���S��\[pCĥ�g���{2��:���Q�Q]2I"/gba����Δо���P}�qC2j���I�HE�e���_�ϳ'7Ż��͠��T�b@3jz�'_"��୮ep;3U@� ��;��o�+�l�]�sI2E�o��1-:�-Y�F�<����x��z�w���Y�����+�_-���0�$�2H�����SE���mk[\��k�Gշf�9�yл5u���' f����b�k�u��^ . �1�ǭ�t��}�Խ1��A���b����Z������x��aYCS��ȟ��IV�/�ml���K����+{��~�]���ѕ���%!�y>4~�T}�\���kZD�,�d������I UX��*a^�q8��}d$)����8e|�c�VYBO�g� �v�|'��t��s H\^�ZT0�G�FJ���gK��l���:��'�I�q��>����95���Z�4>�Lm��(U>�q��X����~8�rq�ā�q�ԉq��jE��bӠ�¿�}�Şd.����x�v��r�������DR����N_eϜ�b�������j/VVM_�X�X~�������8#�F�1}�楩��M�	��B�Yu�ɯ��@�ڢ�r�����s��6Ͷ_&��AV�Vվ�O�ݴ�k`�٤���)��X��A+��0z�Q�0P��^H1H.;�Ś�"����p�oT������2�,�%���3�p�			uI^�|sx����ŕ݌X��7��'��F��� *q��e/ʟu��$�)))�VK*h���Q�?��P���=|E �kf���[GK����&�oR��î�9⹶�|m7*�a; �J�9��n�z��"�3�/c!5�0-�j�c�®1���U�'{�P_|(5{��x�����r|�Q�[��H}R�A�jj���У�Y؋ч�ɴ�����J_E����+�Ȫ{�v�+@9���2@����^\��e�7_U�u�S�f��Alg�����G]Ǥ�4E�������3�{o��M����-���/%E�wVd5jGzƚ�9��~8,f n�*Z�/�`@�<ذ����	��N~{z��(z�}�<��$�z��>��%u���G���D�ywBi��#˳h�ޑ7�*�ɢ���T�%1�4�ш�׷_W�1�E�lQji#F����?M�R�S�ǡsr~<80p[��Usdl��5��	�7o΁�=V����U�®��8@
|���pK�%&�;�cR��j���w��ܷpʪWG��9�/�R�I�]�w��\4) `ғ).��:LTуY;�F���ր��Y�r%�N	7ܑ��D����<٥�P�i�J����R�Nzw��.�1�ҍ��ߜ�=�j���0�����Ӎ��z��7ڞU!��3Ծ�%�4��I���V1��N�SSt�bdL�F�s�װ�
�7@V�l`4���H77p|~���inV��r��jaYY�P�vE:R\p�����7�2�_�jip�U9�@�Q�� ���yʗs��=<1MN�#���e���<���_W}�ǘ��z���K��&�^"��
��;�Bd����JL��$
9M���὆g��p�n����l �)���t�� u����~�#���Y�E��'�%�PMs�S�u���$"b��tB��::�Vۘ��y��Wu��*sU�;��_Q�ٳU8�S���_�3?�:�LQ�w���f��[-�e����p�ˢ?�zs�?�	��kz<�vXR �jW��X����Z�=,--]�,v9�Ϫ������FZi��S�kԕ������i��8x�*�FOhb;o-�荎���f��	��n�7�X�Fu��,])J�)V��i:��{ї1��|�}:��f��$ <a:�͌n��h�Ff�"����~�L����d�+���`���@���T7��|H=7��ֹ��@����`���v��~&��{���Ily�7hSGً�b?K�u*7�js��b��ʷ��LMm�?�WP�'�����`���\�H�Rǟ�|x���69�J�a�E���u:��1��Rq�g}f��xy�F��ӷ������<W�����JJJ P8o#[�D���W:�=]j[H4���˫��
$��������:ӏ����s#�1P��!���/�6��y�X��D��u=��_���IUu�Zf��?�����F��z��X$2ڼ��쨸%b@^��V����*ւ3x���nP��Ou:�
���[�RǨjh��yN��@��Z���߳,��X���c;���*�?�:Ψ������*�������3F$sq���F&�@t�kfM(�*�s_�m0�ݏ�`���s��jȔ^���R�JEm?[����8���7��j�"��6,��!"�6ߊ�.�Gg���_�ڂ������kX� ii�$w�b������"OfpWW���&�}S��Q����,�������H����R9�r!�t�,Q�bH�!:�����K�M��4Īz�e����7������\G;��ҪY�B/�#p����jq!*-�z����΋H8�z3D��Xu���Q�+.޿n��X��
�°v��2hG���2��:6GT�$��n�����	�?;��r?F�1s�>� �Pr��9���V��'n*� �*����B��į�Ƴ~v��I��N��d��}�� ����G�m�L�x�* O����yI��⃃�$q?�1�}dP��F7,�=2��M5��BHKKwTG�,'�X*_*�qŸ��1��ҟ3/�S^޹�BJ���փb�'Rֲ[q�ס�Ii"���IjY�������@��2)g����mR��i���V�3�)F���ƿŢ?����,�8]�V��}����_D��[��n(����
W�\Q56������]�Z���� �*�F��&Ʉ�Hj�A�՚͞�p��>�ȵ�-|�U���>�R����NV�x��MC��ڳ0-~B\��Q3�5�a�3����-���O4��������^�"��g�* 8��{o��:P9������9�'��P0�>��n���7��8�I�[���5���W%vd� ��Y*�]�d�p�ٗ�R$�;=lr�1�c�3��d�&�	St!�@�/J[�#8���N�#��aSX���R�1�4"%$����OM^~��%���(Ak��H�R�=s�,�B��'���U��
RT�}y@�)h+�3�%�G���ְ�Cw�R��H���uy��؟���+�%��F^�y�;���:82ZVB�����{�}�M�q�}����{X��ֽ%�����ǋ�~��C^Z�݃��j<��	L��$��D:eV�}ܶ�5�E J"�I�A�w�GG�	����|��̌ ��:���)R�ݳ*jB`��G��!�<�Yt[2���S�i���`'/x���Ȳ�����Y�6#�FD\H�O�DO��r	=��Ron�J(:���l/^�fXXs?��%�mK��>-�P=aa
��)
/�g\��=��猈��X����)�̥�T_3��{{;�j�C+�-�QD�����*bɘ{W��� ʦ��V,�:�{1ϛ:��`s<!T0�N��{���A���¢W�����2̤g�E�$&���� �;���F���nX�F�'�7�8���y+�{`o��?0��Ŧ7�����uMG|�/2�NǾ/!y������F��Gg�, `4��(e�Ȯ���~g��͛;�U����6��<Ɵl:���T֑���S��H�x�9n�iX��JB�ɵ�E#R����}[! �v�--�ka�,�AJ\@��4$�C�����F����`QN��M���{���}11I��XQ5�Ð�^i W@�����:�����	��?�ݺn�a���rcnsӢ;:v��4����� #u:|�Y�H��I:Ea�7�5�K�|9��?(�2���,1J�J�#sy��,�@;i���g����6a7��<)N��bc��m��|A1׽�=��%0��,����qS�
;f4��:(����Q��=7b�M��M�s��ْ�J�r�g�6�y�=��R�6W}�ً_�זҎ��j�g�rr��{��AY�n#�N��wfj+�xn�1w]G�*�])�%O2饙�Z'�#��RO�_K,�?Ο����Z0yJ�3`�`6a����R���8&S� �T	�1��מ$�؉+	g!"���Az;�{[:��
׊ .�.�djsK�b�O��I<�6w�e�1&-q1�|.������"��E>G�g'�5�^��]�����q.M�mA� 
ԕ�'�O����s���>�2|����0pq���^&��(�����9��T�Qq_�V���ͳZ^�W���(�]����lu_{���T9���mC:��� LP�F>��ԸH��W����RP�i�RJ�^�tD�����o`7��0�Ŷ�`���i+�\٦�Ŗ����DT�"J�#��g�v
��~
FЬ��SO�7���i:z�'�����σn �-Q�L�/�UX�b�M>I�)F�m׎L�@)���N��{��(m�=�7��0������ �����{[���^�!����8����1�u���Z�!�J��׵�w�&�.bfo�:��ڂ����jĕH�x�td_�
�����\C}i`�D�Z
˘#n,��w�|+PE�"W��N�R�>a�o�:c ys�J��	����M��/A/ ���6�p�0JZ�>��H?	a,���hGy��N�c9B����W����>��QSˎ�ᘖ'�k�r�"��b ��Ɍf�E�޷`g�O�*�>z�LN؛RIhOY�f8޼=_%��V�����gw�<l1IÇA���#�=4l T�K�3)x̲�N��x���[�;�� 4w�v��Pg�$���:S��8�֍�ⲴB,�)�_K�Ư ]W��>/߭���aT�l��h{�9��]�|s�5��Զ�������Q�D��a2�}2�{#�8��a���Jwf��t�Xa̵c��X]Yi0x����M􈾰"���L�~��!X=��H���>ث��8���NO׎�iG��ζ�s��lz�~t��hO�q�x�dro�/#��c�|��v,vҋ�t�"�)��~�ˡ�co�~;@3M�"�2�pp]��wg�Z~]�[fs�m@�%S��Α�^� ;�p��ώ�7������H4]����O�*��OL���GKs�zp�PΦ��r_�����ѿ�H���h9����t;�ݏ�5�֚5��?N��Z,,�;�Y����`�A��`Tb��s���P(rr�H^ӹ��'��G���Ҍ����������!��	����|��}��[�Ǽ�ϭ���yr��/��S�g�hٙ���G��,D����x97D�r���9�h�R@����ʶ���D���d*�A���P�	�Ԫ�Ō;�J��NX��Jk��.h��Ѹ��G�4^�[SEWhK�ۨ�E�����Z��C���	jg��% ��46[�����="�(%M";�,��t�{��6�%��ԛ�
�Z�����SIS�� ;1u~n��L������|���v|�qYHmjL����c�yۥ�85�X���Ό�ω_��ƕ]�K����E��b�9B@��It�`�!J�3+�Z�٪���:��vr{=2�[_�}�gjUE&v��7=���`ԯ��Sw���m����5:��2�syQ`�@	.��چ�	�5b�S���|,.���dRn8�t����7T2�"�}lKM"�j�wR8h�ݜ�v��w�f|7������
�v�M� q�!C�ȦT�;G$�͞,�V6�g�xVV�B�����i��k�͡����- �p��=B�Q��mG�>�S�F���8-t=������q������Fjq�B&����=|�X{B��B;��C�(�v��L���]����Px�������R�/�:Bh��N���4��	B���|0`�<���-��p0����C��T���gU�_Y�8�T�[�GM��	� �q�5��R��e3�f�p�r0��K4�Mҝi��B�p(N#�6+���?:3J.���'�m�&x�`p"�`VW%�,n&oຑ&h��2��_v� ���sOXv~a�G�����P:26��[�c��>_��aQ�]��_2��T�`�iS �O�x�����ҥ�Xuf��[�뙢u�k�@@þ�����χ=��)S�Į��N��>z�ZQP$-7}���Hu�hB)v���_]C� �Hi.7��/T.�����7
*��{cWυ;w0�'����<��+�R�Z����+�=�7����Q"|'� )�Y��O�(�2М��3}����-ο{��N]'�=C���)�.H$m}��5U��k�N��G붎�W#:>Ɍ��~_��͸xo/�ģd� k�bu�F��&T��Os�2Q ��r���`тO���������
�6_�2K�bK�=nu�2���S�)�̣�P�N;���q��Tf��f��Ju57=�=�Z*  ���% �:8Hae<;�gt�&�������Ӯ�m��-2�����K�꣭"�Ƅ\�~�=)��N����+
��kt��� g�������_��֥�рI��H����V��t�c[���XQ��{>�r��so���"N{���A�~��`sZ�Gc���9+'��Wq{�p˵��⪤�l٫�?u����Rlp���R-�WC��.���gD�BnĲA!.��8"�ԶP��紜�c�
��k:L=�m2p
v#!�~�Gb�@0pਣ��9m)X����Խ��}Z�'7~eC�XD��N`�f�J�R�bRե�����d[�=�cj�<��sJ-Z p0m���[U��:��>5��Fn(~���s����(b�/�7�Yv�����ʆN�7}dŀ ��'��&��t1���́{��7�O`���ut��ć�ڤ�⯕���$��$��e�[�6Q�C 7v��h#�YR����C�X���J�^��[)'~��`q�閦�����$��qI�� �x��O6�l��ޞ��&����������$$P׭�rT�A���������£tܘ�OTٰ�h]�SQX�h_�k+�ŅJw%g��S��LAFe��j�L��r���;2+��_��������S[?�e�Jkz���z'� hd������?Ƅ	��6Oe�i�uVy����p�KPVZ:������5IB�(5�ٹ��X�]�Q,��O��82YC-�k�R�&�dɲ>�N2X�{��/eq�I��&��b�ٙ�ڮ����d��p/��)��1��Ȏ5���]j���������'pW�#�~�)m'��]s��QLg2$��E[D�Ţc�. ��'4�<CП~�d��� �$0e����%�P���.���������Z�4U�� v�l�P��y��
�H��zr����F���\��HM��������7����F@L^G𗋙���B�q��f���x]��1ѷ�������|*"%�	]�6�	�K�"�G�:n�$.m0F$�ߕ�4�r��'��a�����<ap	��M���B�>����!���n����g��om���6�o��c�=�u��ZХ���vR��m}��:���J�6��z{gG��
/r��IК�C��;�܇G'_��H]z:֑��}�"it�fi���w�)�=c7(K��>���E%�jLU�)j''��Lw:ĭ��`06f��A/����N����V�)���)+�-�$7LoK��>�~a�BWs�=zR����✱i�
Qy����[�u�u�j�U�+��ؘ����j�|?�T�p�}_"��~}���yqY�O5;썍G�_ŷ�Z�y��˥C�"���Љ\���&L�jXeǼ��� Z�e��O%��ً�)���4]M܄ogz��2��*��B^F�Q�GU���f&>y.;�F*nM=��8*j���\b��ܸ�`}�[%��M�K��*�����1m�0m��O��ѓ���;�:A����g9�����d:��G�� r�`�����]�[�4��U�������ħ.=>%*�R|lF�c2k�I1e(�`�Øۡ,O����W7��Kc+��BK�@6|�����c���d���o�Ag����^ǹ�y_=Q�Α�m�)��eC�=��rx��V@��'Y�����=GW���,]�/�Ƙ)�����t]�`;��<_��|��_G�h��B[=�/��8�y�h��ܢ��W�uq��<�R�*�}���c�$+�g�͸V�0�@�N�shDau\�6�8�
�?#fD���0ߋ�6�Rs��H�D΅*�T��G¼4��s���rBZ���ߍ)N�Q�ׇ�ifq�35Z(g(S�K�LT:p�P<��wh���ܨ������҅��,��{�s�������:�|b��YxOJG�l^���Pl'#�}�(�t�J_!n6�-��Қ]�0���Ⱥ`y�x��v�^����ʗm+�.�1b�2����������Q��K��ڋ?�j![?R���ew�/���s�q�,�e��-hZs�s~�*�t-��1�Â���O=�T{�|���7ښ���sA�7U�G�7y9�����:��}�}��8�f��3<j��ZE5���~-N��w�����&��$#s,[�,W�d��9!�/�7݊��&E�a��JM�Mff��V�q��R�X���骩Ň� ��\1O�Ǆ[nI�g��y�L�[��X�Y!��+����Ww�����tT��������u��s�Q��x��u�T��A4H�3�Y�(��=��o%l����_����<%�.nC����w��h"�B����t��۫�dl��\e�f��d�����ܙ�����sZ�=0����[�����|o2>T0�M��;��&�����M��F�<���[�,�7�K��Vo�U�2�|�]����l-֛��BP{�����ׅ��9y����uܺ���6wfz�)n�efw�Ruzmơ�i�Vj�t�` R�jd�~�:a��D>���O	�ͮ�3���Z�c�o�������ش�%ZD�!�y65�(ҙf;�,��r�����J��Ρ"k_^�k���F���u��빋~��s}�M�"q��r��	���M��-ɏTފ��Kb�\��IU!�������O�G�z_�����J�Z�V�!S��	`r8�r�t���&��>���Q�ⵆ1;H7�@��*�w��S?Ǩ�����I"{:����Uu�f1}�R�tM�j=�S3�Fh����yi�RC���K�};Aoܺ<|!����
��N���p)#%�ӰS|�IpפU'�z�;]�I���f�XEo���f���W��!N����$���m�;2q�,�!|o\z_0��k�>��c�tLR�����̠�U���E�xawi`~S����T�Db��X�]�Ӽ	Y��v��L�:wX���mw-���dɱCNQ�� 4�(��h�.�ޠL�W���O���z�+R�u����ǖN.!��"-����"l2�e�5����B��E����ۼ�k��-�G��+ۡ��9�:2+�3Sc��j�*�)�ft?ģq�|Ol�[2�on��߂���x�@�K4<��1��=z�l2~''��
����@�J����cv�o*^��7~��ϻ�8K=RE��z�+(�XN\�@�ȷD�^�]��E�O$�8χ��I���;@D���y�����4������u�e�8�8�xꕯ�u5��\����Z�1��q���\�-��Y`�-eZ2(U}����]$��~lU��ܑ���7�wN�F;�9�p�7L]���<=�l��3�J�8Y��Y%�)_@�v�'Ox�?x�b��{����c����P�t$��]���ꜚ��T\?kI��]�zv�m�E�<��T�P8�dd&�^r�` �χ���2M���6Ui���[�n���R6�e�ܓ�e�Þ�A��'�L	M���$h��m��l�D�_��;Z�q���\ȳ�͍g���A3ߏ|6��A��Oğ3_�;�n��IcT��a�k�:�C�a?���YxkY�����.����Է��*/����P,��p�w�n���TBq*�~�ˤ7��c���C�Zf)�)r�����g����i���{!��a{�Ÿl���E�v͕)��~8����Q6��7��>��j��IO�}�(��u��|�Q��wo�Qu �(��xu��lvi���2���������q/BϕV�O�#�� R-S3C+H�~�U	�X���3QT#��Z�P���������>�"؞h��V����n �R���$�[�����:�����92���yC"M��%�9C9U�rC ��ڹ��a�9�4�lyk� N�qB6W�	�'�E�x޹zMn���P�B�*+�k�ە�P$�(�i���2�>5iN��ԟ�"�t�9U���u�"��r v\�G�(���[cv��w,R\!N'�z]{� #ڸ�n}�V�Q�33��f�����S�.elќo2>`�e�����ə����RTh��Y#3���
 g@���D�l
�55���s�"j��(�t�՟��4�ҵ�����V���e��MIyZ|�SSn��>	H8��2�� �z��sv5^`+����E�}S.]��N8{��Tǖۃ17m&�1��Ѐ��������}����+i�d!t���A�[���?v����[���,�x>�w�x�OOƪ��|t���b@yRrI6�~�c��n�M��- W=��� �ql\y>�T(�X���R��zZUV|zAY֮D{�E-g�*� g%
2_9|�"MB1`�'87ѓ��:���:bn5�Ftճ.%���f���Dd(�m1��^a^S�F���?�a6���i���z���X7-_wo?�2Ά���<@���]����y������W�b@���s��K�+�@U`[�c�D��,P��z��&%L-o�>6Z�8}����Yf�����7|�|`K���Y ��o�1���Qr�9�/b�2<�۲?��_��rQTn��d�o��3��`���ӌ�ƲJdQ �n�(y�؄�?9���V�y8��RiCz>�#�3�����?����%Z�#���8��3*��i
xm�zz�P��� �z�I�j���Wj	-1$*+V~�����4���td�鸺�t����1�V��eX�@��^e�t��@1LX̨[~{�O�q���p�0Bw]�����IoojT�B�ғ��B~�?\�\����q�뫔�C�j���'Q�M���1�;x}��w瓹��e/dEռ�T��i��D�W+w�P����µ��־B���,m�^�McEf>ÏG/����� �LjX�@ؓ���	ݚ~���5����74R"��K�ȕ;ǚ�ɞ�һ:�7܀��ܲ����}�h�S������s��ϱ(;��\R��̉Afi7�(������W��(�D�5<����Ss�0����ׅL��е���q�a�����7&�.T�]z�h �p�o�-�j������D,�7��(W�JΟ�c��q�]��*�z${z���؆���DI!Sۀ�䂣��i~f��7
�K�=�}r�����e�9�P�'%�R�Yke�ZvCg&�4.�-�\����������9x�J�e�Y����q@aV� �+!T[�TX�e+ߜ̯}���2K* �����ȟ�UtO�8��ת��T��Z�{Cwé�F�.�zj�b� �y�����G����v��������H��u�-���/B4��|�4|�G���B�+0C����vQ6����ܗe`Wy���2t��?�"���ѫ��,0�|gz*�^��p�D�`r�nJ88���:�` �T�~lu��L�[B�1�D�!ܪ�聽��������3v�R��+~��4��9�;?�3+]&x����
2j@> 
:�~S 9���rC��n�K�q�	#9�S9n��t�XT0Sm7�%��I�i�<�y|��$��H�)��b���Xh�0�ve���cO�a��g��#&5!�6M����k4��Mo[�$E8{7���AӢҏ��3_h��H���s|@��[u��@�����Pj�K�P��Gi�60�}k,�k`�pϮ~{_�����{�7�U!&6��գ�' ^���%'�&������#9`au���Y���$Ǜq����o��4�?'(�L6^�Q�sa���A����3�d��������[�Y�To�,�`׆&���ũ0�2S~����B�=E �{���>�"|����IOh��,om����|x��l.��uG��t�R9S���N��
i
�%�
K<�D�ߡ����RQJϷ�i���3�=Fv���'��?v�̣�Ŭ��y�\��u{�>�(u���l|�+��P`|hݨ9:���mg��E<l��� ��kM�%',%�ׇ�By^r��-L�%���j�dʅ9�?�7���'����qrC=�+)���J���+���N۰@sE�F�/�<�ƗF�[}�����Y��W78e���`��T��-�,��6�&�󺺻 	eKT����U�ކ��N7.t>N�l+*Y��q�1V��$d靰�;���i/k0�����[l^D���C���۠A�gN�_�F�e��Z�h�a��p�T!�e�	��E�D�UF?��&�B5�XPє2
����8�k��?:�@w%{L��W75�@��q��?��w�\ 4��Jǂ�-yU���#����	���\1��"q���d����2-� [Q_cL�2u{[�t�����Dq�$�q$A2�!��vOO�r�gn�L���������5��������cŃR=�F����?��I�ī4�B�c ^��4�A� Ei���>��)�Қ퐖QQ���W0ƷZ�������M������� f�h[b��m%����w�M�k������}zk�8��[I��k���W�c�r�2l@�F�q��w/8v�������X&�`�@���3q'��9ҍ������bV��l��O��oё܈},qP�f�!�H0��\��ߦ-w�Fh�)��Ҩ\��F0�D �g3.3�.F�O{pyp}�	СʈK�#�~Ы˒s���vr9ic���Q�>פ�f+���9�Ԫ����b��br ���<;<C=�a\#�u��|${�5ɽ��B�AM�.��J���+ufz�\�t�u0�~�"�>��<_m�^j�g�2�ؑ�V �V�4�䗒�k���Ȏ�sPjzZ���%P�ގh�
��j�v����{|/�w۩����I���k�ۄ�����e5  .�s?���7�7����L�`�E�E)�I��r��?2򓥥^���.�\�ξp��x��FO����o0~��ܛ��[1��t�#1�Bؑj5 z����V����2.��e��=���i��.��%ߟ�7.@��RN����(E8�.�+&"r�r�zDg��u�Nl$��,�"L�Ƶ�� �i�k/��1�=2฼�T��O��ڃ��%|z�J9���a�K��7�Ζ�f��gh���7�Mí(��|��A.o���8%��u�EMN^#d�ϣ���=:��6ۅ��6;��p�P�n?���G��S��π��6U�9�P�8h�� ����3&ʧ_��lS��c�*�܍��;�]���	���No<8���3�1��l<�_�z����C������A�69�8[�@����HΪEŪ��ӡ��	�_�Ϭ�>u�sg��[�*@w�v?��*�^������E}"�6md\ɓ��=t�^�B:��=S�gvl�#c}-�^1���@�����W�J���jt�Zq��U��f_��s�画#.�l�V��G*���?UC��z0d��ǖb�
���&����w�H���u����pכ�~�o���	�q]�,�麲��f2�T|����.����غs����-���*����������m���U���*i�Ο���LD��T������ƌᬐ>�>�q7Ap�(�A�P�/����5p|9��o]8��eo7����SK`OI�1S(5��v����1��2���1D�4����� �.�}|:�_c�e�_�H7����DS�� ����2�������'����pՅ=�ٷW(y߼,5}�ܴ#l��cӄ������<+��~k�>�w����[���&�F����'3�����	y��`��&�f`�P	0D��?4�]
۸��eV=��uWOψ��4cu��X���~�NeނB��h`����� A��ϩ��j*i���x);�;�G�=��OD=P���uk�{�����Ï�;B� $��n���ҍ�ޖ)���G����o�@-[�A�r�����A�X{=%}����1����ܧ�%~~����3ݞ�B�V@� ��Y9��Z���[��y�#Ȩ����N��Z�4�s�"�n�T,�J���6����| %�3?���3��6$'����[�?29���B;1�&�j�C\�Ř�eu���w	;�6uJW(�}t�Do�`��آ�@}mN�BSq#���h�W��������N���/�\Ɋ���&}�,
J�F�5�-���9e�ۃ�/%%�ڴ����u������r�dM��/��m�ɭ�o�c���N�Ų9���+s+� ��{�Z��e��	)������p�v6��񁘦i{�?�XaIy�||||�!Atӯ *�vR�{Un��Fb�j���%������ /*�@+��Q��An�V&��؟���MT��&��"dk���XE�����{�a��/�����.�Z��TؠS��,ڔUb����ӜN��2�ku�:ES�̗׭5.+jOӕ%+�9,����3O4fOv������n]X�������U�w{���nt2ڬ�9	�0"@X�b��Ւ
~��W����6�!���3��O�ه��v�{�k�8����8�5����:�^99\G~�r㦮����S�2$�W7d�� ?�{�ӈ��?�O�H���5��,��!�*��ھ>*b!�((�t+
�4H��t���) !���]C����C�4CJ�P߽�}�7k�d-�{��g�o�i�,)-��ӄm�6V�Gr��ű�1�\ץ����ˆ��t�	9\.-� |2�����/J��?Q�d�#�����F��%��PJI,]<<&�x��[��-�r�������<��T!)�/M,u���	&Su	�6�QQII	f���6{�Nɉ�ބS!!������WU������9sٙ	K�kT�b�#˻��?{��o���Ԝ�ڌ���2?�
�	U�W������å��=��:�����sLn L�['����c��ʋ�x��"t�W�$CG�1����K�t��d��ڋ�ل��\�c�t�YL򠨐\�G�e�V��� Ҥ7�����T�ׯ_�l�h��#�ֺř��#���w��]c�� ��wV�����b^�xKP�j��pX$�����a	X�-�&{�uttȫ������
�{�U�.��Ω�B.�:W?��� )�U�;�LH�����n������"�D.o,�Ǻ�K��b��x����m�������}�a4r���e�8���Q�3_����#Li�c���=�GA��ʤ�Ä���D������g��8y� T�mVy��A7k�,�h�H�@�\��8��-�O���:%�iJ�KY���?Rz�\R�|�������o���A�F^OO#�?l��l�?'���SW�"�B�����{kj��8?�Қ���>	$K8�0�ak�AW�?T�(���@��
שj��53�<����"�����ic*:�˘h7����5ȌX��tu#��q�g� ��[c�v�kGB�э�+ Ϯ�� `7�m (7dTPR�\ޡeb��t�c���V��m��~�
�j�[�������������/�C|-��F�{0�
hl�B���I7͝�o�J�G���Փ�<�t�:�d���d�C��F���E�W�с3`� ���e"��R��


FM�w����\��&4�{� ������(��	G�9��7Y�L�9X��+�;ou�)Z�g��	��c����b|<P2��f����r��랍]�ȃc�q\2l�����4~PE	�!���[�>���:U�g��ʩU�8��־���yю�N]9�)��%%�bS��B��L�bؖ�O�f6�#�5��]A����  ��_
m%8�?V�Ee�R�K�&s@�_����Zk�b��Y��e���|�� ���%Ă�Ab�Y�k��(��"���z��66#X�.�I�j�D����A�V�t;/]e��jf 2��W�O�X1���g4����BC�?9X�L���_��7�A���;j��}�V��hpQ�,��4���aؘ�����JL�7񦚈W/�|�19��p��W�G��E�se�sE�z/bSJ�I�UrdH5ૻ"�����������!UJK���Y�>��$%�dʒ��!Zsω��Yc!}q�F�&�4�2�i��PI}�G�l�� �)����.W�Gݙa�)�$���U�E<�gv�|�k����x�����k6㷽^�c�,1ZIz@��u�����?���I�(��M�ҍ�q0&XA�|'�9lrA�{A�S�ESf��u�rʞ٦k�����9/(h:$K;���4�v|�Ǧ�� j�n��j�~pϮ�v�Nx(��P�NjǴ����7���dH���ތc���eXD���a���%`>ǈ&g�\�LI�V�\E�N($�}K%�_�ve����/��Y�}�1p�w3䤸(�N��qW��^��j��o�p̌���R�8_�[� ���!\��Y�x6F9��Ny���Ck��ё2mq��m�����0���눿��n�װ�����7&{e[#��}m\!�}|�l|��0��8�ɘ��)߾}�<�oZ�9����Om� `a-�H'���h	��ڰ�w�b[�宅�)T��P<����-6��x���o����pJ�C�S�5u�=Z�1��Y�cS�b)~A��I�lR2Q�t��(L�s�1�n]}x> ��{R#���Nq���_	�N���Iå���-�R� ���@��4�ZmQ���o��]�^���L������gP�	�I�������g�N��4��f�ډ�F�YhK��‿��|aE�5	�W��[�L>-g��1p1v����@���,@:��$�ϡ���i<��N*@����Xn{����WyUb^�%��'�k����T�����w���q�1e.(SӃ��>�V#��m�FX� ����( ��ץ�����k�3���0�l�+y��N��Ǽ!RB���2$yt��&W�cQ�KRv@��P�t婤����d����!��f�q+Y�/�f�j�?�[a�r�|ߢ����e_7��;�Ⱥ�����l���zx��>��c��<�����,���Q��X��x���[�P�f�L�f*�ƈ�Hjo�p�Ou�??�m).�@�ڻ�ʥ9�i�Ke�쉧�,���OKG�oVU	�6��2����@[�9� ��M4�WR1
ݺ��㟔E���䑪�7�&��.��ifw��^sK&؃:�v���F�f��5G��8t�7���$�(d�w�\EBİ��8N��`}�U��&����]�o	�~6�9R�a)�B�1���6@�;���K�\�;h�'D!�ҏS�\�y�Vm\��r� >���N��BY߫��V<��e6,ُ�t���bc�O�]pDiY��Sѥ�`uBL��9s'��z���|�W�Z��dE S-\����`.z7'q���$T�n�������kre�S�C�,���a"��|NmIrc� 7�v���QF�J���+�4�L��~)]ŗ��$;��9�qX��ɤ٢#�r�� 8���$�\Y@�x�� � x�����6�����j�IJ������S)��o��4&؂��;�����-D���,�OF�[x�dd���)4��α��$X� �@<�Dv��,3��V{��nػ�`��V��ɉj�\��s�\ik�r��n�L<��<���NI0���%_���~i�KC�3۸1�ы�����l��Lށ��Y�U��Ԙh����ޤ�tr��&�:'Sg��1�-��Ҝ0�MKή�7��t����d��X_1=����9��[h�a|�MYW	�S"�2Dn/�Ǜ9�2�+��2��ItD�����%�a�9�u����p�I�y3J�0�<��*�.N�|�9i��}��Y{Ԅ�@�yZ��:X�Y��n��e�-�z3*
�fxg�����:��0��	���yq�l����(ꍏ'� �p�$��2�g-�Ӄ[�km��0��$+6��)?�;u��b�"��?+�D��D��K~6y�B�Y��ȑ�W���cW�pm�`��>c�A��7EQ����-���f�����$��6Q�`
�� �H;y23(by�RLǈ}M�}����4%b��O�N͙E9��e#�%N>�e25`!a�Y��[��x���:�b
���5܍��|��=�"�[!^��{$�����	���zҨ�W���#����wR��(�X6mֲU�����{����~�P�1�r��{�����I$P�(�8���n@����2���9���T��O� s�m7���Erp������Bӈ�ΰ�&e��!�C �m�R�%��7'�Ʋ!T,k���v� �3�¤����ӏ<jLآ�[.�o�A~M��	�0R��8x�&� �f�P�k,��Ǖ~�X+��(�x�w��j�2�,{ӊ/����	�]�O�<��fШV�i Ɨj^0Z�5��a!�w�"��G]j�������O���BT�z;
�R�;8dU%����ZX�KBG�b��
�ȭ&�s���|��;D�櫤�/:�R.`��oQ��"
 h��>/3���~[_qg��Lz���E6pYI��(��$���kvF]R���=�!
�Y�uhΧ�����ۧF�8�C=u�S��Aۙ��)�~ݒ�3jW�γ�"箸�.����թM��l'���dn$�A�6�7��x�,��ߔx�c�Wn�esJǆ�q�Q�U84k�)0�����5�z��xy٢� u�&yו
�O:/�U2����)4\�Q:A�qJ�����
%c�$lt��<�v��
Q�{�����sBJ�._���N1�ϙL}��|�S�{Kv�K�O��;o��L�S��ce�W�v=�*�WZ�x���0�e�����u/���]ƍgf3Tl��q��JГ"������ |+�J�����G=�D�J��]Ж����rQ�N���Ǫ�1��\"?�2�۷s5����`�(���C�<\�s����Gtk�G6W	��S�މ��/1^�zn�T�9{�OJ�; ��播�����[%;�J~%�H�������_�8�?���O/[���/Č���};����yd;Dݺ|m�V��s_}Q/ J�$o���FL����v�u��Hߦ�6=��͞xr�q�i�%��^w���qg-� *�J��#m�R��
]�RZm5/u��ƍa�"��\�69��so �v��-�z#���FCArb���ˡ�A2�u�v�Y�lʫ)��q��.��t\jH(��9��B��̒��Fp!�ʗ��>���y�)i�IՉ�=�J�(jW�<k��y�x~�C�A o�#FUS�i���H�w&[m%^Otp: )1���=6(yS��>�SO�*4�f;v�Xa<�
�j%wu  (|����!�/�mY��av�b��-4���a�E?��	�3�V 3�+|s=���o��S����8�y>��u��?��'2�+��;?c0����>�*�ǝo��M���$4-1�_�e�·���W��c"ް�*4�5�Ù��x*>�F�x���C�?�9�c�k �|�2��s�t���-^_3U���"������`K��'Y1Sr�󛞌�7ӒΩ���a��-$���T<�'C�Y,7uH{Ow(Z}%���L��u���d��s%�%���k�7/��ci4M���C�&?��k�D�V�}"�'�^Ae,b|�n��o���;p_>8:�\$��d�H�Bߐ��Ҝ/�=unD���V9�x��qu<.���l0��/!��TQN���*�Tn�#�ψ#d-aɜ(�N�K���N	�~|�����*R<"�N�OW�q�~s1/�\���(f�qX�&��X�=���O��ݝ��K�"'.�K���G��7wt�Cm��u�ׄvl��YXXX��7����nQ`y�$�05���� �ɑ��:��U�䱙Gl^������5�d�X�7�V�&�3 �uW�b/�^�6J�G��.Jp��G�cL��@<ϴ��o�ב{��S���ף}���U�M�����zg.u%��=�f ĩV�Q";T�12."T�o.k|���Kc-�"ԭ=0���*"�!G��+�ǯxx�K�^{�e�k{$�8~=������������ܕ��)K�&�z��+o�\(�}���,��S3灁�A�޼���8��jc����j�3λ���3� G���9�]21Ͳ�KpX���E� �q�:��Lҿ!:a�>.ǠDB��1.�aP yv����ʀ�y�~l�]f���������O������`uJ��f��^���˻	�/O"��}��ƻ�Qi��V�ջ�.�68{�%�8��-*�"+�\�,+:`�vS���8�dN�(ބIv�)LI��9���'^���~����@�� �Аgs��t{N��x�{�U�]��5_@�����f�$��E������R�z�-��Q���֥�ƺ�f�;�Ā�In�B=W�#͛��rpm�����ȇ'�dp�Ro��5�v��z�P�5G<��^|a6�W��׺�~���E>�Y4��1U� p��VeU�bY6���
��to��iU��
��s�����@_�9�I�9!LE�$)ve>��&v����˨���p*	�$�� ��x-�n+�@��݊���Y�Vx����/���}��Q�'nO�l�7��jG.�h�)?5��V"��ƣ�|2�x�����_p�N�ȓ���ol���~�3Q�#�2yp���:CN�% EN����7E&��+��f�fP�r�Y�+���_��"C.��T�T�+̡�/?�2�Bk���S�פ��pr�h�:6y�ytt����H�����eء����D�ź*�3��_%�+!����4�aA�o�&�
c}<x~q�qP��p���}�/�~YfbTi�m���~���qR���,ߵ.n�����[��ѱD�]4��)�ٞ<N()Y�[i�yc�P,#�k���C��cr�nI��� Z�*�N�C���;ȡ+�緈ZZ�UY֜���
��!\�R�����P���.cS�~?*0Vn2��_9�LDp3��'��H�QGw����7�H�6���)|���7L��ll45�mqQ)��gdy(��H��N�Fp���&�R��!�7$n��H@��X�L�S֔���!7�Oo������!�?�o�o�c3�������d��3����a��`?}���e��>�=66x���H�p�?{�HK�����l��������Љ�ZX8�{̢�U�������S33���gQp��d�G��z�ផ�ryv�#�z|�OP�^'�s��o��;m{ݘS��.c8���ɢ'��mć0��hNB,��U2��*^!W�d����):U��ED�,!h��}��.ԡFZ��T#�ñݏRV��L��u�Y�yëJr8cZ�V�e�45���B���*��S�9wc�L����"a4թ�t����p:������5;#�߽".�|qw�UZ#�&iYvS�.����l)m{��Y������_�b�^Φ.�L��r꾃�ѿtΊ���]�R%ا�CGO�)�姨+�)+g�uFа��`��m��Lq8�w#��I$b��Չ;%���+�{ꃛF�w�a���J�����/����X��Ka�������R�11��'t#���(g��� ����?+�b�D��������/��#Ww�ɞ��1}ݯ����@q�֚0��L��oI���N���EF�U���b��l�b{��zm�!d�w�Y9��Q�*��09���턜�z���?��e���Ӱ�{�x��w�f�7��l�ě\5�n\*e��\�VC=t�ed|drA?-S |ٰT42�@��7������|�ω���2Fv�d�uL�捂�g��dvaAd��G�.}�l`��+	���vi5=�5½|���B�է,m��td����^�%�/S�ꨕ�w�%�u�@Q9�D��@^�Y�N�)��x&{��Ң�U6�1��}�3Ipd$^�5�Ϊeo�1��h5���INJJJh9Zi!��s����;��]�p�4"v��<@���[����z+�8auf�.���j�9�;ZK��Iy�^5�c��t7�zh3��;� 2U�+���}꣐��=�;�б�,���)7F���j|�H�Q�q��\�̾b�y0dҺ��h����}|�$�`,������b/���(���(��4�Yr>���'טkvK��+gn���ǝSN]�h����^Y����.�q˗G��\�$%%�^���p$��TY��5���_�GY6��X�<=���{���O"�� �51����lш���r��7jrI� d4�x2�FX�Iq�[��$}�)L��x~+��,�o��Q�O�t(���������`��Y�϶�t����m|�9'&�4��Th�3�g6�
�z�br��*g,!6������^y�=��c�/XU�kh�sc�cYZ^��{��#z%G��.���ԓ�Dn��zG'ώ�*�8�]�4��B�=��jF�o�6���EqL��,���\�OINV%,|Nd�b�;���D��R��i�A�֭Ӵ�x�)~m��k
8������J�~��������G�2þg�v�.�s�J�jp?��־dЬ�3��ͷ/PX�2��wٹ�t&��o�4�A�#$k�F�)(�W�Ŧ�t��Wl�;Hֿu\�����v,�Ȅ�Z�ڐ���Ͻ��������w��(]��#	a�΢9��nL�g�,O�R
�U~��^|k�^Y����wcvn��Z����Z���R�V��q�ꧬ|�?Ku���zz��1�}��`?e�|��:NK���N�gAX�cwm�_�jNmQ�"9�i��z<���,3>�鯬98��"9��;8�x���ĕ3H�۟^���XASM�*6z�;ȍD<���&ώ.��v�K�F|6���nF1�C�A�}�A�+���7�p����T��UIX�6��.Q��.��a�g����r8��.+��nR�1�t��F|J*ۻ�sq��1<c�L"lW���PW��677ˬ�:�"F)� +�&��P��4E��k�+��u�J�$#T���U�K24�e cQ�v���U�]��7����!��Rj���� R����P�9P:GM����Ɨ�}	]�,V�2<����V[�g'7�6�7�j��ؗ�g�1�+:�H�v��+&!�L�~����=�ͤ�Q�r��g̗��j��������E9n��Z�P����8!���=��t4�_^u���"��TK�iU)ZsPB��d�@	�$�\F�KX��f[�"?�S�阱����T��:�3��z��|أ��	�h�������m�+���y@Ġ�Ln�%�����YP[[�U�&'�
��}Bdu���n�V�tj�XʥU��h��6d���,���8�u��Yz��Nu%�9,��cϢ�v�P�<�]�;3�6K��?�N�O���G=_!�6"o
S?�:B�Y��K��qq�0BR���c�� '��ӳ"�$��R� ��N��HKZ5L�K)!v,��J:�K�V5����*d�.�ua�8��|���CC-���B��������
��-� &wY��*\ǳE��~o"��ǰvw���O����w�k�g�-Kv��&9p�]���&����:�f�]Ч\��v\0����⋩�I�1��Մboԝ����ۋ�A�f�>Mɟ��1��GDFf$8P.��6V=Rj �?�fv{�*��7E�S��7<�>���%���I�_;�����-��@&Ջ����՚��V���a��O����6qo���Xq�ԫ�RW�|8Z��e~�NBpP�T���	#?�������e*��������TJ�Nv
S+ ��a�4�*�=��촯�l�Y� [�4��j|�/x�r��_:���ȸ}ÿ$�lѧ%�^� &���pS�G�t!Ŕ��C����@�B���A}1"��-+�g���Jpx���jOA�\�/]�|X|Z5L}p�.�|>v�H�O��X���	����ş�C��hT�j��0~���m[QG3:�g��k���N�V�wV�H;Q�^�X�ˡ-��O2YM�o"�ꁦ��07����S�B*ji�T%#��(���roDڬ���侫�A����8|qqdv�a����H��%1F�B���J_�Q��L���Ys����T^/��y��-�)�
�qy��2�S�%u�k2J0�����$�pO�6��sd���N��Y�!8hҺJ�����hE/X7���T������D�W.@�B;��&~��/kB$�,ȃ���mN!Cp����bӱw����]�
�L0J�b�uR�+����-�t�����u��"a3&�˝�"�2�1����uUn�1���-�!|U�[(�-�L܃/x���w����?�Yes��
��_�d�q�h�ڳ�q���e͓�<i3r���.��k�;W�_5F�����\�w�^�`�}�qE��,�R-՗����g�ǵ�X��J<%g�+�^�l��oVОx�����N�}����4�h�Z
�D�mo��ֳ��k�0q$厖����䢪D�&|�*=$����$�U[�|����n�Y��nv�i?N,&���R٢-n=Zì'y� ~:���$�ls�n��PA�����@�]�� �~�@xK
��r�6���褴�B�>�Sԍ������W$���$Q�m�O����B��%	��9�T\�3{�5;ē�bj�u�8TR�K���o�a��U��S���G�Ʀ �w�@ހ����c	���o�&��,����ܭE�LI�K}�x�x|����I�OIc�Wʫ�YUޘ]-��M�T-��-�r�Y6�����x}�+��dn�:>eo?� �E�ʸ9��*p����T���PX�����ܣ�=��	�j��l³G��c�uEȪ�|�����}{���o���@o�SiơvFm4k��jO�OO�c^:�D0�e477g�!��q���K)�Ԏm��My��j:��l��h�5��f�k&tN�|Vf�$�V��nǠ��ѓS-�՞[�褣��`_M9{� ���
`l0�f�����d���9>�2��$E^��s,�l1�?B5}UZ�\�^b��>��[����k�;���u�4��3�sϤ���>aau;q6��ck��V�E��W:l�e��X���ly}�T �I���G Ϩ��|�`o��a���W^�q=a1���O����8,�2�7o�X�:��+R[NR�v��ұ��Q{���a�&�Xl
��_&�Y�I���ٙ)a��yi3�`�Tp�ʠI�u���r�ol��(�,\��d���*F��v��d&���a4V�q��EA���A�h�i��ā���
w�������F���D%C�n< ��)���y�\$�P��^X���
8�x���>.{�	��ìS�V6[z\��X.�R��Q����)q�r�놃. 'R���֭�H��K�#���ꂂqC~�D��]��`r�#۱ҍ�Ý��5|����S�e�F%Tg&�$)X�:���fj���M���Ig�8��d��� K,�.uĵ�oU���k]c~������2)�f;بx�;^s3�,,�˴��3ȳ^��`c��qYC ��Q��֋{	8*Nf���wm�.�� ӑ�Z�hw��`K�/�37��d�"g{1+����ͪ�j�p����g�<C���}��\ER��5�+l�;�z��0�׈3�e�\�8UK Cs�Tj��S����-I3W�N��o޳6Lw߭��n��ݕa��_�6)���;g���b���)���l�B��\�B��_~���v�b
6��{��jI��`��r��$��@6Lf×G�Sؓ�3�ձ�v��qyvR�V
�*�ļʹl2}a�/C:gTB�ʳ���TM�<�z9R5�إh)��FM������@#%&�W?)��T��J@�&��x��6���k�7��`���t?*����N���� �,$-Rӕ�x�Y�7擔6b'	QQ���q��ޤ[��+J�f�>�LMJ��7�������+G	
 n�YEg8���j4D$�ҪǼC²�3A͆���uX��1�,�V`g��Sg��P�|	�E A@�[�5���a$�����Sžj�7r��[H�$�v����
XE���m7w��� ;N�֕xq"!��܆�z����Ϫ5#y�����4���� �G����2�ֺ���JO�j��"L����|���½��ŝջ#.E
����0 ���\��j�>4�@*��y��g:>'���d�W��m{�w�s�ԛl|���H�u��<�9`ᴕ�ZӾ�HT����aJ��vNbib��(� 	"�߄s�l��� �c�Y���闳�L�;�(��f�(T*l8q�x��g`���LT��\�!�׻��+((��D�A��^�����))��-��о��7��E�:7�;���P�7d7�ش��������^m`M��L.��`
�UGc�.?[��HU�'|���J�7^����C

H�[�Ei�
c�t�Q�*��(*�嫼������f\�����&B,փ?�7<rr���|��4�̶s�yI��0'���0!q��[˱Y%q�wW"�բ�a�!�BL.��^R�!��x����7
l_I�)7ۓ ��{,�ux��Uk�1��t�x3*']G�P���S%"}gy06�
�
p���<����FO�.G��������>4���I�w���ci/�E����07�p<��[�I���=1� Z^n��Vs���+�,7L~<�k�9�<���E�"�d43�4���q���W�Q�^����޵;2�ٰ%ʱLv
d����DC���s LC���
5�p̷���k�y>�{�n.ݯ��k�<�y}3�|����g���t��R����҅������MVɂ>��2��EAuV��}�.Q�2��\}�@��b�$ ao�e�@b1�o�G�F�����2s�=�qMB@�⫹<%�}{����]�^�D����[�@� %�4B��C;XH��o�WK��vE�n�"���dŤo�G�؍�鏗��d�c�Z�jHٱ@��'���GgRWt�W���=��O���9D(i��ٰ�J��h��w25�){���KFdu����_���	���Z:u�e�3�����ܒj�lT�7)D٨FvZ�[�x3�W�c�Dh�R��x|��r}����;���^�RI�jZ��������~B���v���Y�����&��{7�c�T�����|����w~C�5yR��T��M�]�\O�+�S����������žTY���˙ ��6������$0\8�#�t�y~��㞠�3�f�NDw	�t<���Tc�:B3�2�on!�}���H-�9>�� �-4S���X9	9�I��0ޜmW��J''�ZS��,��|��q�!��� ���ޘuP&����I�5����Xs5O��~�nd*c����8e��S���w�ư�k~�n!`ܳk��v��<�#�4�v}"?[.sɏ*!x�<hi��`�H M�(ߘk")T)�o�/}����&ù�����zU���^��o�Y��#�F�F��O2��=`���*�_ʛ��]�<&'��;j��. jS��C�tz�����t�h�6�a��/k�t�,�U�Ӹ�D����$]\�N��m���oV�眒�ⰰ���AFi��JCkP�f�7 ߞ}q1�� �T�յ޼�`>���|o����`Ô��$[����8ظw��1��
ߣ�&�/k�_�Ҕ�C
��Ў�R[k)�[�	�Ր�I����X�И�6���<�}�w,#�;�q��z���T����vG�
�T"���D�����6��j��<�"���hP����k����^=���;XS�0�o3�Ϸgҭ}��NA�P�{��r��������?Ȁn���5���PV���x$YbO�����c����
��ޤW�̬ 2��u+'7�%�
�S~��/����71Q Ji��Q�g�}�?X9�
v�=x��v�I�Y1lz���ai#�3\�V椅"��i�Bخz�(�)+H���$[tm�u����.}��h��7xO:r��e�m���rNK���SJ�eED��-�YkDB'��0�����v��z^�o+))Vxd�	 }��u����*�݇6[]]E�;^@�Y����1�^&��D 4�1�UC�t�[�SԬ�~շ������&�rO8�Y��?���צ��ԡ��,|{�O���?4^U�����fQ��e=�X���,w��:�zpU�����#�_m���N(d��Q�*l�)��L>�w7*$$��P�uf�d,eä�5G��qq�) k����=`s\���x	>ܿ2\��]��h�s��|��F�t"_+3 y���*���c.�	�V���u$��&zYjǣy�=�г ��|^��ǝT"�{�-\�b[����H$ *�777��qڮD�W���'�u6���>�լ96e�6$_h����߿����Lk�dd�*c@��X�y�nݺ�8�MD^QQ�^��h,iﬦ��N���,�G��v��8�AB�RJ��Ʌc�Ō��<�T�}X]��u��jfHDkC6���hU[�+K7@�@��i��dd��6sݿ�^(---d!��dW�[�4[�Ϯ���'9c�ӓC@.���˫������{�,'���fA�k�N�a������Հ�)�n����{L���`'9s��ԏώ�;� ǯ�[�E3�s8o�ˤ�_��r�9�Rб���!�kT<x�d�_�-�	v?(��$B���c�,���`[Yx�i�s-�>��H��B�c��'�<g��,`pD����$5ł��'Ǉ˭��B'�;o��m��� /1����e�05u�6�U\~|�@���K�U�S��a>����s��"-բ�Vl�Řu;�m����6�y�j�ބS�ˡm*�t����rVf��Xvvv+��P� <C2tr�#�J�� 8S ��vNN�a�=}��ꨒx���bD1�G�b8-SFFF��	8'��m38���5�M\�u�73
G�å��SR��<161a�����Ύ����?��Ossr`�v4Am:�>  �u�L<i7|+��mo��.�]"�~e�J�;=';�Eĕ���4�"�Ѱ��.}��Ԥ*L�S���S߻��K�r!��!� �R�.���L����1�F!����צ�� K�Ml*12|�E8����\2�Z�n��U����R�����k��E!�������>@��� �gȍVGʅK���v�� ��B}�gJF0��T�I��8l5��/(��ʋM�N<�E��/�!d��㫝�YN)����C�����G�������#����|H�EP�n��O�t� �y�r���w���G������~�ip����)cO_�7a��p@�G�n��H�zhՖw�W�dt��1�m�}*�z-�л�oٮ�0��W��R�}뢼�-:c`�4HI�߹ ݏ�S�X�}� �X�~w �LIX||�l��.�3�-�[2�тg�d�ƕ���v���Y?6�B�da�!��tTk �e��^�[e����}`�*�����<K��kԩ����n����j*�8�zxu
�1����w���\�O3T>|@S�D/	���b��v{�J���_<Z��ݻ���SIu=F=����<o`L�����h�7<f�û�s}�����ܫ������d�M�/p��ڱ�����������A|D�T��:�(��KE%����c��p�l�zhR��{�
�n@o�@_�����-e�
��5;����H�8Ȓ�A|��%_����.�+4/���{�V�����5��&�;�Ik_�K�޺����A����~��eٴ��x4�t�k�b#Bm�������f��,�?g�l��꠶��,.�<�%�6��_t���o���$*+�/�"W@8���XG!Wт?Tf'i 5	+�p��,Л��Zz�� �#�,7e���'1�/	�K4���\���/�%^� J����4-~
�a��$�J]��K���)�/B�j���a�2Ia��J3]l���v|���E��n	���
�65gT��R�n���YA�X�&gk[�aU��v�lBXX��S��#�޻�8ᴎ����o^���g�DoU	D]&"C+���+�X�Q쪲|X:6���͘@t�V�4n֚��%ͅh�6�t�m���"͐��sa�tc��5�,��|~�Z$g���9�`���]j���5l�+̂��u�`�2�[�ט������8.�Yl��t�)��w�1��j^�b_�ÂJ.<L3�0���Q�������D�;H�V�(�=3�k���4���g�@�Ʈ}r�p���7��:`;eն$���B�S�!����n��!��a�X1r	#��v�4"�?�&s�4�j�꠆&������-�?���_6,gV(Wm�R+q�S')���+'r�L���� �*�[��%yYV��i�J�o��@�z.�w�9?�p��_UG��Wp�;P:�M!�)b�J#��~-�4;�-����*�/~:��k�e���*Jp3|%��sf������V��g!��	���F�QI'�-��F�ᕓ�j 
fP�?s)��aq�F��_Z�Ӎ�T����'<t��u�+jʖ?�ֺ�[]󕎐��<0��<�歾�X��i��\�f��3�xO�ioQfߞ��0���	9���#9�o��e�u�Kw��)6_��UسY��u��d[	�� ��j�H�ؽ��a�h�C��z�Mc��0��=��.N�gV��* �@��kT�3��=0.J)y{��'��F�r�6VUM-`��e�fi�������*1��4��G�1r�Hǲj0[����"t�T��۔�𹂎��r�Ɂ������p���_�X��y&g�0"����C��c?#9��]\�1.���>-x�59���l���ݒ�+�#Y���7g�v�f7�%D���|9��&�ͳ�=W��ښr;��X3f%:;[ҥz���ڗ ���H}�Rk�E��r�����98��Vm�+F����ҁ�(]��R�W��R�(���E�6azc[�&�=����@v{Ip-��!��!@N�h$�UW^��oJ�V�6�,g���y4&�����>�	#9C�"��b�D���=B���(��&�3�����ǝh������m�ćP0�[,�s�4N��|>Ȍ����HwY ��<ŕf*��r]�I�4�ˡ�x�a�~�	F����r>������"Ξ�ѵ�e�F�Zn��D�;0m-|���eg&�����A�kv�����1Wi/�������}�^�*K�Q�U��H�a��C�%5�Jok)��ֵ�;�=O�:8?�1��26�\n��3FRJD%�����B(�FW=�j[��B�� )ɨ`dd�w���\>XH� tٲ�݀O)�^4����(ۓ�^��8��<�=�<Ӹ,#W�s���A�8Z@�ى�� �Uת�v������3��'<��'�����TUc�N� pPH�"5]ă�~�����Z��0�x��F�����Vs9yeZ��#=9�y[dz�s�vHZ�7b@,�0�Zo�GF��U�o�Ef���>`ym+��[&��B'IVLd�Y��g���L�9��u<G� V(c�-��U"8'�E����I�/�����&������,_�=R�!S���@�ՅG����9	�䨖gת���eW����4ߖz���X�
%0�o¤�
�6&&�F�T۶�ɵ�?+��GL�a��e���O}� ��L��ϟ?�iy����������a���j��:S�rT�k_�ٿ�X?TMp�"&$�O޺��@Z�I�B��u÷W}�m;3J�� �Tb��qr�o�o���C%o�/�#�!�T�vt�,��	����[ 2BR��w�� w�!�S���=��-��x�MO!���*�A-��"��X�����g�r����KbqHa�ƚN��Af���*�Fdy�Ob�����͹�p ��W5B¢p11ج�%���zݽ�(����M���i�� ��EdL[���>�LB�9���Q21tɣ������?�)�����"+#�C���#[B���J���$+�d�B��Ce{��{��p���������Ox�_㺞����%L2{���Q+�/oe{������g��%:�I��>_�/�2-/.�J��D��}A�P�@��-�
DB�9/N�n.�&jpW��A�����z�B��5��@dٴ��.g&����YW���O���:�k2Mۣb�k�O�]&?C���|⽤�m>+$����s�F��"����S*-��>+�+qH�;pܠX��G�=a�`��H��}ҍ�"z�Ϗ�������|�d�����3ƚ��΂i\�����������	��w�*�����"�O}��ج|���Vg��5r������T��;�����ȉk�`�3]�~hbz�wu{g~=ñ��JN��N�Z�!����o����� ��������=�!�-�z��x71����aULX��,�ӗY��Z:�im�n'��Y ���"`�4;;�M���b�kHYYY^��#����,Gj2Ra�p{o��:���jl�(�/��Gq�'�}�l=R�a>��ʌ���)�8���o`� ��x>��3�juk?<��<#��8�a�50{����vk�bY4�@a���`P��~_�*;�[`W�]nCxs;��X�x�va_�c>ctz@�-����:[�w�0�2��00��H*ݲ���bJ&�&�*S�V�4 V~Na�o����\� C���\��/�����a�2�ĕ��� �*�7GQ�J�"�:��������E�1�ʅ�u��W�[t3欏dv���j�х��=Jh[����վ3���p
�E+x�<װ�@����&�,�>�����<�*�9`n��� ��-AA-A�s8�U�ik���%Fz��q�b���[;���J0�����7�p���������4`�tB ��Q�A���@���Y�O7�/߇6� י���=�I��f�ǼD<lſ<}�8��tU`Xϡ��3��UJJ�3�ev�qx}�y��~@�"�[C�WW���� ev�4=p�Xe�N�bh�~b��G�s:z�B�,S��b�9m�Tm�r-���z�%�x�=F;E@��O�zb��V�+����s ���ϣ�P`$���\LFJ?�H<��`�ң QXBs�Lz�E����}��!����q���ϝ�����,�l`�qz�q=���qH�Bp�;W͒��F���t^t�-?Yo��0��XD�^�N�,�f#C}[�L���ɭ0�o�V~��<�<��a�y�� vWvN�c�מ�C�Ik&ֈ���`�VIÜ?O ���l����{���D!��P�)�=��	�v�SC֚(�b���ᮉ�9�5����&��Mb[��������P�̂�Lz��AM�B&��/87!>�=�� 9�y�5;��|o]��7��5���"Y9_:T�8!���LA��� E�(� ���C0�����	�i�Q<�>qY|������V�����$�2��u�q�@$֦��	t�-g+�_%�h}A���̑�8n^����d��硸J�r,D���P��ù���fg��?th�����KM���Do؋�)�0��6Ő���5��y�B���~-r����:�Ϋ�N�6���T$���R)G��v���d���S5BW�q�1'�ө�����w+��,�wi�î����'�b�+��lzlF�$M.��K����e�����_g}���Fύ�B)��
!��Y�<�ߒ��
?؅o���A	�/���l�|�[�"��W*Q���
/d2��;1U��Yέ�]�=M�f����#�Qz&"��[��17$BZ�ʲ���r��BG6è{����t����"ց��xڄ����՟Յ�
��^�\���g3��-�i)��"��.N�!�g�9������vW�Ӕ"���_� l��������XJh�4��-s\�K��z����4M��Ϲ]����Jo��*�ś�
(2R�����<�%
#d����]����뼪)�oF���+���zR���OK�CI�����j\��~h�p"I�^��jio[���sM댋l�k<����e�=˸����鄪�:;�No�W���s��m�#ƃ��Yj3J�)�����dHl��z�u�Z�3h8�7 ����8��=L��
	��Z?��5�鱈/U�w~cK�R%%f��8u%w���:�.7�����UN�z�+�r����-6�Sn���0�R:{CJ���1�p���2�z�����I=R�H����Gr+�S��aO'w����ON�cS�΀�o���N�l�_��t��e�~��+�&ë��:�L��>Y�)��/�|�d}�M9�D>X���M\#F�i�hY齡,Ów��ev��]4��'oEۖA�{��cA�VV|�ǩ[��g{_GI���*v����Y��M�1W�[���Υ3�=���2�f"Vx՜��\���� C�1xsd$����������M�[2&Bme���P�ld� )�r���C��s�o~@�@j}�����q 1�Ǽ��0�_�r�(ի;�0��g��N+��$B���L��|j �T�˿Q�ѺҀ���S�{�lٟ��+���jc��"9��'�H���^�a8�M����ٹ9�Y1��߽�S3�̌��5Uݻ
*rCW�ߚK������?L���x?j"�!sG�c�uGw�2����w�e�V�b��|fJq$RǏ�˘�<b.��l�\�,/��_g��S��zU)�������Z�ܷgY�+�x��G@C���I;�$�3Y�Z��ڨ�a�5B���D�'Ӿ�癶ju<û�J�:h����`�*7�\�~ޱ��������PV[�w�'Y�w�v���J���;���g _�<�3�8zp����mKz��/��ٝf>�,~�ok�i�R�{dᖓ.6*�G�oEp���cޝ�)	Ģ���T���TB�L_΅�_־�u�(I����-�^�+qn�$�hVi���cd�7R�#��[���'=��ai�b�%�U��~����(�3��hͳ�ҔO��`)"�Σ(3О�S�WįH@��Cȝ��jdl[܌�������]�3�������M<�~�b��OT��w0�\�B6"v��T'�IOV�Mm~/u�a������m"=���Ԩ�Q���d�D�R@~�ku�:��?�xN(ׁ�,��ғ|v�m~�F�5`O*��uKƤ ��l(x�P�V]W7Cg�˃�ub.] ���"w�y�Z���fTAEҮ�ˁڪh(��h*���e��S[M��T��l�i�u�\T���5-.K�-�:36������8	�t���w@�� �}JW��9��SV�r&�a��ye���n�WIz���v��S|�N3 c
G/<uSz��B�ҁ(�|��IA��ʚM��a���z7M��#;-���V�r�[�D�����A{Oׅ�,��j��h��Vn�t*q�ׁ��cn�KٺA(Z_�`;/�~^�����������W�b�~��ZjwO��W�+�bq�B��L����&V�Va�Ǔ�We�J���3~8�Q?��x	ߵ�����7>(qj[���d�,v_~9}�τ]~�D�0�v�ѕP�n�l����/�G�ϖ^�r�aC�#�:��ٞ�E��?bDu��l8:���$�f��-!�s�,�����aBtt;8;;�y�(�n���$9����������k��u���!wk��4w�$ux�R�0��C��4K��%��c�%���Ș,���/D�|����dO�#��y��+H2�W,�e��B�W�36����Q��F ���[����b̮�sC ���мN���e"r��Q���WT��ԙ�z3�����L?��ˬ��_���1-�Ztʺ1�f�5�����GL���#���<6���C<N�]j�P��)�G3ї��2�� ˬd&����zL��NOtm����;�;�X�}�g���j�E�ZTO��ﲔsB��ܔ����?�B�8��#�h:Pq����b	햳��ۜ-���m�huo�v�ie�wX(*y�e&`G��w��&Rr,�0R��`�����L��:��v��s�@��k 8�:88(?;I����f���u�����  9�n�&�1�d�����^v��D6��M}�%�&;G��)[��2�z��z-S*�	n^u�RȎ��"��@22���	� ���)'���Lh� 11��45� �j�,�93?ϟx��o-`�1`�~}L�FJF���DL��Y�%=�ff[���-���F����N����r�6�yxW<,�z�J�:��T:|�V�M wblX���\K ��T|��p�4J]	`���7����݆�����DFD ���ӯ����W�H�ae �ee^ �\h�km�1�ѕ��/n����K�9x�o��x�%��
�񥮭c�9����Aw�Z�$�N��l~�TQ��Ȕ��@oW�|��/<��a�H÷��%ϊ1U�mjRq�z-THc�{#,f��JJJ<�
Znz���HU8e2<]�C/��͈`��K=O�OzN��R��.����U$0dc=��lN�:��={&?5b?�bt�v���W� �Q;�7�����?�q�_�b�6��@�o��z��Ib�e��U����(��]����
�u�������*�Z:��"q� � �9���TO�8��Y��Xʷ3%N?o�GJ��Dw�n!
P�څ�7@]t��T�(K��ΰ��(yæ^F����?t���}��5{�
=[���\2P,;�v�r���z����N�Y9����ɓ�!�y�ZCKk6�ed�~�1g �e[�m�elY%,������[�;���.4�6:�p��!���w M���=���;4��"o
�s���-'uT��?&q��9(�Z�?�䕏9cR��g�Ie��֚����AZ�{��c�1|�kYl�Y��8|*���D��ї{���y������9�Od�nӼ���dX�����5i`c��&8,�`lS!+�-���b28̼"-�w	�H��o�.j+��`�*('X��L��u�������3���0�@Rf)=�M�����^rQ�9t�[B��X��!r���ϽC�7�31{� ����{�n'�\b���L�y�.�����T�*�f-֟}��'��];b�ya�#�=���yQȚo��y����**)$�O�]�*�펏��%��m�J��ws1�	aY���fE�����h��q�����X��L��.�s
�x�h�(�W��,����~��aǅ�\`����V�9���S� �w!�*霿��p,��JV��O`/���.��O�o�C*�y��w$ͨ�\|5��&��~h�)�Ce�[�c@,�q떲��ّ �t&{{�xl�g��8��͊^� 9��f�x9�y^��4g;�%�% ��S2} OEYݩ�Y�L�g�]Y{��7g�sF;��[Zx1����ފ���gB�gvf�a��V1�����Mp�+6�AU5�/���"�3�fm��(!;��&^�,��Z���f�K�����������A���6�5� jd�z�T��K�d��B��)��!x;��j��.�ٱ��8+��bCy�'�P����ٝ�S�U���aΪ�K�	-��q)KD'/�� �D�� 
��\�g��G����Ml\�)׼���������� .B-@y�A��?�V�.V7F"U�)��F�0F�ʘ��ˈ�Tl'���V���D�,W�T��
�ǀz�H��)�I=�I���.>�'ru.�:�˪��W����r�y#����d���w�B��X���	>?6 ����U���Gd��і���)6�`	+�T�[Ұm���,�n���墓����h�u���Di��}�������E�h���T}����آ=�<i5 �����r�"n 	QF<OD�Xe� q�t���ۡ�^�̀��>��q�����ωS5��ru@Lk
2br_
��q��	hO���0b�I	ߢ�z��U��##�L"��Y�Z�y�ށx���o�{#O��j�1'��p�b4PVY��C g����Eh����wS�R R{8�Y�)����s.�w`S�~��r�l\�I(�uQ�����=��*���S~ĉ�d��]9�},ਗ��|j�?��2oe�y��W2jkG��׿��jI쟋4j��Ѷ�l�f��<�rL�}�c'A��k�*=i���Zg����1�c��Et�B�xGcm�����_�z>�����X��P���;0`!B�؄�VꚚ�p`�}���E��*���*�uB2���Gm<H&��a瘝de{#8*T ���">��zWbs��`�z�JWR���E%Kp�'�{FQ���3�r9���_���)\8 �tr�,�?m�8X�D����-c�Ȝ �F��Rd�4�y3�3J�	��@`ݕoed�1���*�dK~6}�5�Im�>��3�%�����s�F�5q�wh�}����g�<�*++��6m�4�I��ϐaUL��K/����u�iSm�^�NK��Uj���Y�~���pҀ�v�1B�Uu%�v�r}�cH�Q��@�K ����/Nk!ߌ<�nQ�KJ1Y��@g�982a�'B�Tn1&>3~�E�{���V"�jڍ!Z���IO6w���)8$w�)��9e���T�:��	Ł  �wfx��'m��H�x�;ʴ���b�t����)3�[L��b/��,,�<R�����f��`%:��`wB++E�����e����«��x�퉒ף'F�דn��_r��7,;W��R��I���9�p�RK�UU��I*}�+,���3�t�f���J\�o�����}��p�
�a�,��yW�����w�=q�Ny��+�������v^w1�!}b"q�����%Zú.�5�����NCA%6��U�/v��E�����'4����;(ȕb�?�Qc��/_L���V�`D��n�r0�� �����m��,ws,����`��R���ի�����e�U�����y���̠�i�����>���V�r��/:��aVB� r:_(8����8�y`@�BZ֛(��/�m����xxT�o��pLzo�g�����̨F7f�NFX���7�����g��-ʰ9����h�v3?��z���|�`���	ۄ��(�ͬo)�}~��ou�d�	*n���_=�<��1��y3��W�c����@�4J���k�?�㯜�Α���>��6P`Qd9hp��*�A�w&�ܠHb'����RZE��S��j�O�*�����pv��sX�y�8o��Eg5Y,\"��'T\�0_��а�u�$��]3�%�+�g��9@Q�g���A'1��*�X�Y��4[�>��#ȕ(ޚNb��}譌�[�'2Zk�DzzN��Y��MH��?�8���e����M� ��½��It�-@�h�.\����?�k�N�|��QF�_�,����C� �����fx9s�-U*��h�3 �L��3�,ޱ:�cu9\�D~��	����]�z�b�_܈{�ϴU=R	�-�,�Ɛ�W�
�-���UZ�EɛJ�n���SH���P�{ҩ]]\v�'� ���Gu���? k|�e�}.��ا"!dC�(d���|�V?��`L��4=�S�L��z!�b�<�F���0g��'�a���Z>К�\�i{]/�S@�%�@��D�l�v�ۮ��k2\���ˏ9�IД�\���e�N,�����E�!����wXXi��z�0��NS���w[˩H5�\��P����ɒ�4��Fj���(�)`	�хo���7+^)�j�q!�l��#u���T1	�1�{vL������BH�Ӊe���r^�l�%zw�c�)ʈ8����3Կb�5���`g�����c1�Ghr7(8C^���DCQ���h�&RK�o��\.�M�F*��P����q�� �":ь�:{yE�k�R;w��T�BN���|��o�K����w��*�M9=I��P랤�q�e����8Յ���� �'VT�V��|���m���C�$(5WH��:�+6���5����:����7Cq�p�;%5]��eu������a��v^�k��(k�K���0�.:�%.��{�^^��<�?�;�(��z�2�)E�3ݙ�c�o4�bt�'zlL׆G��ʤd��n�h��}��Z�QOgvuY7]�;0��
I,{�l��w�s�0ǻ��6!FmB`p�����*����v� 2�g�p�τ��v>���^4�K~\6��Mf�����3�Cy88h*BR"ZvjPM��&f�������Z��O|�S��P-c��P�>p���r%k���A���	���Aɇ{S+�5��U��`?�l���WR+;���u�w���C��X3{=��5��p�]�����T����[59��W�Adt4Th˗��S�6�����⽿u6q�r��(��ɒx��zF�>C��͇>�~|��Gva��P���pq�]X��QK�%<oؾ�5�d�&��YG�O�ݐ�줺Ȉ�3!D�;����YU��쪻�qI��r��-_rz���n��H[5�\O
=ձ���R,*Q�cM)��-x�5R3A%��r6V7u�hފ�b�b���� ,Tc%O�3�0���=�x���oԅ�y��@�ؓ�fv���^����V��SI�OzP���aH���k�Ū#�&׻�U7��!�w�2�� Z�MI��T�h힎$����NX�+)�9|5�U�[U':6Pk�Խ�Yu�7�;t%��O�kbx> �)��#�����;���{kY���⁉�o��D�A��,V�*��2�ku��%��]�h��mˬ�)�rC3�鼿K�v��)�>�|��׮�����>K���Lo�<{ȪQ�C���2#4�9�ڣV'�A�����ah���ǀ���^ס޻p�B\��bML���1o��-���a�;�;��֗�Dֺ��N�Rw~-"ߒP��<v����h���8�R�r���E�;�N��>��iZ��T��wN?��w���c.���ٌ2+T�ߓ.���X��:�.���J>�9+q��B�p����"0�F�d2�;s�9S�>��.�h7�?�H�$ͮ�p����g.A�x-�Y$���`u��f�F,��XJBM8;��M�s���ֻcM�)�HY����������.T���{vʻ^^U���1g��"j*h�[��h!��U]���;�����������#�����+_cc�*E=`*��c���'ۥQ�T+v�#ʱ�(�E[���<�����S$�>Ć�ͻ��%��}�j�~��%���Ӛ<؜Z@�X�D�n���1���]��\��,�Xhcq�� ���h)��ai##P���no�S-t��qƭ��rx�*��Jm��=�El̆'��J K�7�^��������l�LD���%�Fh�s����lBǻ�6<���������oB�՜��ϕ�]p��u��Iiw���X���=���+�@� q(8�t��̏����U��ij�yR�����\v"������B�+��٩]�
bO~�]-5�W��K��ڬ;��;u�sr6VVH+D� ���~*�����wH�K;Eٲѝ�9�(}^��g	q�:؄RNzc�6� aN���P��@}��>At��!|��.Z��o�}}���B��S��)�>1�2���	]<�tL���V�n�F�������Sח��(7	1�Q]��<�)T����o!��͢�ػ� �U�k_ϸ��9���1so
�CbB$%-x&sb{*5Wgwi�}�������J���!g��y���ꮞ���֝���<F�|?�ɥ1]��Mu�`C�pxv&�E�]rz��tVfRO ��qgWW���`�]r�HubG� �[t����SI��5^����7��u�e]0߸����X����	������BH�d�A�&�'k:v����6��B�-,��P{�32�.\�03;�fe�s��7��Or��H��ܢΞ�,5~����f��H�.��m|f,3P!$>�el��-����Sd�WN�(^@	������$1/ys��������[l�S
�b�f�}��2Y]B�%R���^Cؤ��:f���LJ
B5�u�t�A��C��Dq8j��N��b3�PR�w(�>��u���ԯ�Q��=KD�����<ۄb���obUu��j�.����´ֵh��kGO���',-��z/xGo�F�q�������b�z�f���L��WF҈>����DHrÌ>�n
�\�"Q7����1��>�7la�����d.�a��^��tIH��x�G��V�����eG�?��e����3S2����Md/	nt�E>��|n���?�4w	3�6��F}ԟ�Z�-G*��R�N�����CX�3u�i�`��d��|2Г53ە����JҍL��QUU�B�����KO�n�X\�v83U����ח��6��;�iiD�B:9��	��U<��p����	oJ`;�u�jQ���[���~�mиw�=��Y��)HgR���ֹ0�j�K
N!d�FM�	��_�K�^ M�D�Hf"舢.u�4X�&{.�ѯ�79�i��掿���rc�K<�Pp�:�|�� �ŝ�@{ߏ��5Y�M�kw�AkJy��<���^�����p����|��[Ӧȵ�[� ��v�?��B���4�h*�j�?�,��9������P���e�%T�{}�����GKf����!�Tm[ՙ��m��r`�U�(���4O�J�Q�ۙ�[�C��P�����b���}w��+��<y8����w�⺫9$Jn�篣(���S|����;9_��s�y
U����:���6 =~��^�޾v�S�=M|	�h��*n)�Z��5v9^�ﺙ�K�C\1�>4mţ� G�o����{�X��S�D���m�7t��U:����Qe�L&�/�*��.��>w.} <آ/��v��W�O|�'1<����G��� �����Ҁ�`����&�;�)����ڋ��������h�R=h����Js��JO ���E��e��3F��?��v3��U�����pC��[�*_��D�O�wۉKh�E���"i�_,YCE-��^az�T�h���Q��eT�"��6^@��sor�c��@��'�1��쏇�W.�(��/j�x�$?��}�V��9X�2&����jv�o1ﺑH$�G�S���^Ȣ:Q])��/�a�|�⑈� _��� E���*�i��<���M�+v$N�{u�<Bt��48I����n�@;@�I  �E9:E+���,�(_,���5�����HO�����ϓ%^bQ�KK��
���CT���C�{u���m/!�^�R�h Eh��\_�?Y�����s�<G~\��2���-�]��z���)@�Aiii��_C����ō������o��>6�<����8�D7��V"d�.��kc�3(���U������z∫h��[��P��P aL�y�� U�o�tU��˖;Lј{��+,�6�p��6�����������򙁯/ٖ߁����8��^u��?�^���[Z��"���m�{�x�$���p�H��b)��Q��A7`OP��e��d���Q�v��o ���[&��A���+�gQ��y�D�G���
|�(�o�K�NļI]C�bgj�4��ֶv%��:p��x����a���ۭ�v���q�:���'��${,4B�.��?T�ڟ���;���ݟ��[|usf�Rl��";?� �p�^h���V���i�`/Y��호��|�S9�(6��ϝ���*��
ȱ)��`���7�y��������l��b��^��ӯ�g�V
��C�yh[T���\Q{|G�]�<����<���.3Yp�$"�G16t6������Qr"��є[-ŏ�'	�i�q�@M�~��-K_v_��E&<]��6���<�@tdDD��fDDtgfn���صޝ򿔚�@�fs��qs{��[j	\,��ߑ�7+�S8{�>|]�9D���
Sg�X$�e�^
C���=��s2���
���N�bI��:�O����W�� � W��7��{Ac��I]vx��4*���'���Ipk�e?e�\P����JL�E��ܟ��65�B��96 @hv�ڵ�ƹ텤�UwY��� H�̬Z��m��'Ђjl��ӫW�b;ө�C��ml;nu9!>{c3��<�N:�rrP��Y�E�.�'w�Z���A� ���H{>�:���ּ�Yڎ��\��T6(�/֓y\:� ��,ߩ�E/��'��nw�?�vtqq����OV���Sc�����j�3��+}��(�A��"��H�R���Ƃ��0�z�X�+ �wp�0=�_���`� ��E�2����}�o�|�!嚹��BE�P˄y;]��N�>��.	R}�zݾjo]2K�����@�0b����"�6[�!��o)�*e�e��Z��mI�aߋ���n��aw=v))����!E@]�s4�z��}1	��ceS�8�K�R콿sL;{�ꍚ��Z;�S��M���۝U>��(N�մ��0D�%|���ahz������Fɇ�\&##өr͓��`~I.�z7tR��{�m�TK��tL��s�/�[PP�b*	Y�9"jv��xP��]��T��L`�T�r�y��9B�*�<R���g��@w^�bB{��SX�|��U%"��:�a��ں��q�5�O(� ��t+��]�wsg�(�7����E�b��'^�1 ���`��0+�+Deq̰`vd�D,?s$%v1`�C]�P3��`���躛+;�
Z��m�]�� ��.]5�X$v3x
�f\)H_�yU�,ɋ��o������2��f���hp,eT�xVb�^>ߡ�����D�7;T���G��s�.�"L�����_�I^"��@w�@���R(���O�c��hm}Ü��2�X������^dԏ�(�Ϊ����D�R��G�n~����YH]���Wd�c�F�!=&���r٨�n���L��$�E:�!_6�'��qOp��ODT���p��u����KLO:_g�"4>}}}���_i��9�`V��? � m��.~�F�P��v���h�?�����!f6ڠ��P=s6�u�eg�H�K���}8`]j�%i����aI�.<��$Յ��Er�&l� ���e���W咥jl��F[5\A�4m6�X\Ϧ��=���S�I����l���<ݲ�*�]����S��dg�P�U@o��F���x�NbF�G;݇�dӝ�l�0�Zlʸ0�XK��T�G����JIF�� �}���n�@����0�0�hɒ�eJ$af�����E�"���;��R��b��a[���,���[F�U ��Ӓ��[N�D�g���w$�&�w����~z��m��0]\��Cx�^���!`��Ȫ�R�Q��P��xC?�I{,�(������%�F�4���"P���Y�(J��������] d�\���mFkk���g�s����e�`<�#C��u���|a�$j`��I�;mU��	���%?��i�qý�B2�������>���{>�j�+;�v6'ͬ�̬¯aj��K�{�C�����G�z��9c�sz��tR$�Ɣ����ܦzVZL��,Ӧ�Z�g���&ɠ��'������N����Nv�#S�.�ZP�����2�������j��Uk�N�P�D�L�BX߱���ή�}�9Z�C|��p�o��T��m���h�2v:#�b�zM:�
��*�kS_nn��ϕ����|��I�?z�^��iw~s܍��]��zz�6F$�^�W���������;�%y��*��U�Jm�V�Ӈ���M�W-���(��/����<?�ǳ�O?��Gw�QM�M�e�OP�F�s�q��%Jҗ���]\0r�;aؓNf|�!�AAA�ۓ�%ƍ���ŝ.Uh(��1`6�@���ٲ�}:�6�1�%����n�F�7���Jɪ<�bM� �������^;͂��m٣�v�`+�I�4��/�}O�6���n��i����%�̴�{[g���j�����w�M�Ug7m����
���Y���7�ܺ7���+�7��7�ݒ��I
�~k���Io9����\����X�)"5`��0���]�]C�7�N�ul�肐ڔ�'&���
	I3a������R ���Ɏx�*��9�W�И����'��/&m�P����:iMp]�����4j�Qt_�Z��9�
��3Ԅ�a��S\&I�o�Sۡ˹А8�Y)y�zh���<��f3�ÇϽ(C�(��e�1a+�o[5/�����1�	JPpa�0�����D�<�9��D�R���1�]�q��A�V���s��,�\�$S�<=noTt-��/��[��3��B��d���s[5�"#�o����)L׽�2D�ա#�|�S
�-�R��#k�(�!�N����gTxyUq��9���;�oO{ҭ��$A���d��0��}vYM#�+�ڽ�{muw��ʭ޾~�켼;6��sH$���y_A����ଜ��w56C�.}j��Z�5ka �.	X�,�a�.P��6��Y;:_���ŭ��-+�J�g���J�ī�f��ҁ�Aے�B�3�vRCKW�
��-���4␰��3tʮє�dJP^}�>n��`����_1}�+��
e�(�M۩l~|����u�5j7�p�,tL�%�9,�	���⽖Z9�_�$%5����ɹg�n�*�g� /���w�JcK������<�����CZ��[��b�>N M��x�nܹ8+���/v��ʫ���F,�^�� ��cϜ��*�A['S��֚v��|�� T���?��9Tf��\ǹ�~F==}���*�.�8@L�ڙ��2�]��˚3%b}տj9Y�_���%��y�hO�4AG��=4��ϭ�,�?������~�5�`��q�F������c�`�}�:��s�{"�k����xl�^z��2��!z��zP�f����Ay�>alY�<ٕ�]7B�r������CϵCP�~Q��Ss"�;& z����O��\K��M�\-nF�v�6��J]έi�A!u�����F�UyYB�1�Y��.�����P8:�`�G�}`�	�f/��_i[t��s�ٴ[>Y���	�� ��uɒ�����rPx�R1dh�h���婏��ξ�4���}%�6�Y��{���gfg�W��~��6M����#/��\l�U
�T��n?�w�ۓ��o����&���t��p3��k�/h�y M���������%�c3g��`jǠ��u��C����-����Bwj8>1��v1Z�^zpX1^1�.�'CPfq&_��=��3�5~��~��b�WJ&��<ֿۓ��Z�4�����n��GA���Ÿc/��\�ը)�N��~�l�3����-J�M#����Sn*���6�o/N�`��2Uy��P�bb(J�zSQ�2&;[N_�{i�}���i�Q�kw��>��==3�O�2U&��>�>��' ���%�[�j;3Zu����wԩ�˯7-�:�a>���%��2�z4؆s���������?s(������H��A����ý26vg-L�_�����������q�5�0,h3�����iY����?�gZ�%_�.����R�[a�&]�@��3�>s�ʤ���ͤ��*�?|#���ڼ�#7�]N:�Xk��11��$}��t+��TZ��g&o�{�e:r]�;a��]���� )�"�v�?��^O�{�x䢯�Wr-ᘤ�S^�M:�l�ӊ{��<?�0xb��f�ǥ}�L��K{�+"��ν�y�m P[��6�h�A}԰�&��0�/y>84�ު�z�j�#����-6�+Wh%[�.��?+�j�z�.^h[��6�'ok���z��-�*��%?C�<���XS�\]_�S����ש�;D��<޸���<���C@Ƈ^ر����>�*�.&[W�{�E�oy��W�vT�_9󸿓hFӈ{+ii�y(�r<$L|�r�(-�������0Z��9>�6���ћ�#��]ö�]"֤�ڂB��}��Mڣ�K[�
�^{��9Co8�2�:k>���r���=��wf��ݫ9�5��}����*�����OB813��b����dʋ�2hƓp�����װ����@���$���@ww��{LD�x�1#��]J"vix37)����s���P�N��03��;&D{>��r��If���`���,��6��󔠹cW�Swݪ�%�����/#��cC�{l#s'�?{ !-.��'��y��g����v��]:vt�*r��d���S�����仉h6�J�Hb��$:et>����ȘH~��x@������u���RbJ:z�kaD�EJ;�n��LU6�}#�[�eͅV߻��#)���MT��%����k�C�q�0[�l�lrgr�X)Rd�����OfnL�C�Ю����'�V�X���Hf~�+5����ݿR�6��plog_����vxp�؉㚩�_f���#UA'�8�+Q+��L�+8����ֻ�͕�|��t��s��j7ۆ�eWKkY�^�Go�%�U�,�Ƨ��E�_QN՜$H:1��_/���'CB�'�8!���b��]����Ȩ�'�/�Gk�$��w_Oo|\�V{�m������Ì�?�f!��U�f�U��R���p0��KZ*��üu��%'n��u@���9UB�2��c�-��A�Ж�]u5�C٣[k+�Q��%��*:S�3^�v��I3ݩ~�?mV*�*��_v��/_���2�^su�������+g�/�
q�b���J��|�j���:l��X��4t�WmJM�K�Q`www.�p2>��0���u���jd�Aى�����Z�ɦz��M��`(��n8T�^����p�XDf�:Y5¹�0�TP$�D�y�{���ܪ�1p�-��,}_�>���L��_���	�
6&���������@T�1ol	
�P(��U��EW�n*;���l��8������5�t�6w4�:T���!���ަ�%~p��Ю�Ҏ�-i\V�e�3�������\O���'�ő�D�Njj��X�� ����\�_=�5aD����#�b�<]t-��?Qi[O@#߭�2.�缮�
�.o���<��SN7a�X���dI��D������B�(X����fՒw"����ɠj�<��;�����ӳ�]���4fz���C��Y��������t9;����W�Ӟ��=�S�h]t�Xo����m���'yJo�v�]�S^x������\j�zp[|Ջ^G�����nv�ޗ�� yN*]�T��<���C���򊉄�}��	���YN`[�}ZU�6�B���QWos7�y�xd�(z�y!��=�o���
n4.�*�I�{�2�g	��}L2�a��jJe�p���y�~2�q���.��q`H���ԝ�C���'�v�f��<i��N��ޮb$����k��w��(k̯�I���#;�C��o��yL%B���oN,)�k�d��k͊�����agƤt�C�}AI���Y0g���������l�Χng����A�T���a��o�M��XS�^���+'1¬��L����y,��}�a�i`����ca͎[�=�t��s6�4�`�6\��R	�6��`��E� �W��^}������z�ݜ��Gl2J��=�J�ʯ��|��)�W��}^�?H�X����M ������r�qs@o�ۍ�Gg�!m�Q6e"�xcU��z�\O׾�u�)뗽���u����f��8*IL*���ۆ,��kDV�}9=7<=ʸ���>��Fte0�`���Ƹ�6=�ホY@��G��'?��ﭼ-�eV���r�a��P6�v�d�;?�?3֔A#�\�gJS����y-0�]�+�C���?y���yI������|Ծ���;a�s�����i��ժW_Reb��s&�{��M�|T����k�vP8�9��]�xR�4N��x���R�'�0��6sa�� �I$3Y��fC��8��4@O�SO����~siD�ˏe��{����/"VYQ�[J�|���:Rk-6~�G+!�I�s���#4�H�R�K4����$���_���|�I�-ł�e@@�t�s5�/x�mQ�y&����#�!+�U��iaw[�N$�Q2w�\�ZV��p�1 �ڦ/?j�p��'X"��N���[����>����{�*��}�xDiRB��PA�D�tw7"-� ��{�Hwwl�κA|y�q�:g�1���ϡc��{͹f\�k��֣DE��f�3�eRp��l��nM�OAzx��P_ʓ�+������|���� �E�f�ա{�&5���Q�5p�dP)���ݽ��R���,�*ׁj(�@�}��c�sq.�zx�>f8��8[�ᢾځ��oV�fR=^�C���4�7��B��?�m��V�7Sor -,�*H��	��{���P+*�Q��Z8�_�E�����>+*���H�	�ߦxJ��O�]Y��7� &���{�D2��N��&��;��ٳ�/�"FC����>Ɵ�N�'�$N]u�xZ~�q[ߖ���(mS�ӕ���F��Lh��٠Uwö~����ڒ���V.���?���̹؟�r�� �N��W(����4w�����A�TE#�}�|����qO���n�k(�濂r����$g�K%�����P�[)n�t��8;��!q�3�&�A�j^3������*��˾�݊-bV�I���d��r�(G�q�X��З*m!��J�P���{vP��-�P]��j�d��dH����I#z�P<��[;��J�ޥ�u��j|�y�+\q�Ml�_o�?>�P-��*�ai�8�����="9?@��$�mI���R4!�b�4���VۇV]��{�O/���:f����)����T�d�8��[����*M��O(7���2m��mt9�h�R�D�� 9q
 |>�xd�C<6!Qv#΃J�|�i#Մ}'��k@ۼ������ǰa�|'�*J��L7F��|k���;Ʌ;^4=�蠖��������I�&�����&'Z��ҥ�|)$�z��U~ h�=ܮ\�8�r~s���5ߖ����W�x+]oA��,��.ETs%(��O�9���H�)�
�-�۹%��1%�rBZch_�{͕8�Yˡ���-��3� ��s���� �mo��._�Ů �� ��݅�R�G�����ғR�(D��(z���>���%Q��X&F�8��#�|�� I�����G�}����U���][��R�i7Y4��?�T�%n�s�z`%��_%I����p��6
jm�/�����
�ՙ�mDH*�2�y{R��QP�`��=��(�9+�1��^d��u\s���/p�׫�0�*n�6������C��g�+���й���@d�a��@���:-�>q�~1>O�n�vm�ɚ`��@�:��Tv��7:Q>��&B�~�����S&Ꮋ�1������OC�xr.diՊ�O ҕ�� l���!.��+�|�8xԸ�zl��3���ťϧ"L 'T����̡21c�� �=��0o����[wvϖ`RW:��� �G���4�Eq������K��˨>�)5�����F�n�ҽR53燖����]^���M�w�#����zH�-O>A��m� z<N�T��4�L|�T�]T�)]R��MC����q^^��~8(+�ֹ����u�D�k.�����l�'��>"��@N�o��"�d�-ǖqlW�2�A���n���h�^�!Ʌ݅X%���{1�R������FO�wv_
��5l���o7�]qZ�	�4�s��`o�TI��U��w�|5�*w^>61����>���	���C��^�9��Jw+����d�t�u�"8ˠ\�`��@Vf�Չ��^�"ǽ��w�`�#FFϝt2���K��|���l�r[�Z8��;��ڮ���s���4�0�١��W� daD�W[jU M������:����NB��Zg����k/������'Gpb]����z1�� �����u���=@k<m��kC�d�A#Yv�κ��O��Vsa^�ɒ�����_E�� �㪖�)
�E�\��R��a/`Im�̛T�e-�X�KUrj�G$жg��M<�4�#���Egz�J�KOLL<���*��d����xĭ�80�u��T	��e=�Y�ό�/�"Lr>��%ut����y���yl�w]�ߔ]�K�Qq"�1ҝx��E�={�{Л$��^e��^'ͦ�T��Y#�/���FW�cG�+��]�zI��2�,�@݀D��Kw�w�w�L��<�ЏWo�&��SY�9�d���R�D��Ǡ��q�:�7�������������B:���`���6��Q�`I_٧�7�ˑ9,#Kj=l,[Lj���E�wP.�g�����`�M�N�!��l�xضg2����@�"�g��A�:�"(%M�M+W(���cM�(x�⹇��ꤔ�ƥd<��e��r{ƺ~������s�
j�nv��	ٽ���sƺEF0w���,�W���*l�ل�/h.�����ʎ6[��gC����@ߑ��6�j�U!�`�����ׁw�
y�g�~���'�B���GOL�1<?!�_BVeu�=4��7���ZDA�yD��Ź^����gӮ �޼�js��s��d�ˑ���:w���|ҭ�r���`v�I9�]8���r�FV��������QL�>�P�G�h��,�c�u��{(6K�{/}���O����>]uZV��^,�UQ�}�����5t�1*�(��5q3_V��D.��;��Y6�4�Ԙ�ta?��Xf�:d�W���>�4�|�~C�Fg�3�4��ڼ=S�Ł�4Vץ�Q��:.���z*����!��~���.����}P��t5k��$�
]��3���8_I*�.��"��ѿl�K/F�>ܾ-��9����JwI������oee���DZo~���92�pKū0��ن�v${qc��[>'��nC�@���ݱ��l{�a�k܄�<d�W�r�=�wz�G��8�x9	#�����G�^+)E�2����dE�zd��[	�
4'���W��+�(2�^��>��t���M	�T��n�4:�Դ�ļ�#��O���	w6N�չ��_i��ƋNSo�#z��e:^�g��-ah�_G�=�-wZ�\r���:��S�]!ϊb</r+��Iѱ)��K��h�/�姊w��_��"aru+��Bկ���9�\�ey>3����%��re�.A�蕷-Ж����U��u����0�K��B����W=l/&��yv�u��N��}&�p�٠aw�kB��h:B
�%��Hz�og0�mm+*�>�:jE[��L�&F��Q3<X@��M�Sg�U�n��t�p%:��r��i=ZV��?�=�C���E{�Ɖ:��xQލ[T����5� -�u�'��4��!T
��\�����M8�w��?�1y6���Xn�_0#ͳ�k?P���]��|��DD1���t|�5w���"��_n}r^�G����F���B=��Z�t�4�d�g<�t1�זw`)J��N���MT�ろ����$�Z�u('��A+*���3�~J�:��G��{����*F���0��'>�{�������F��l�ѥ����֫]>D\ }�D���2�F0R��`��E$��̱���ɸ\[b7m����8��.�r�m���\Nt�o�we���P�ؽ1��;��1/糩��r�bw=��ֆ_R�/�o/�*�Ď_��f���=##Y���#�Uf8�5t�:�F�U��]F���˩K4�u�6��Ҁ�j����ȿm5��RC��e)��t�+���	2�!�R��"��s���B��$n#���b:��?�]�}dr~�	�k�p�Z��")�&= �}��cATis�\�6N�p�M�#�Q��-1��1��T��c��D�S9 �~��Z���[n����-�D�t�.�rT�\.��8W�3�?�x���GZOP���=�hn�3�kW&N�Wx�mf��|��̰L��s��,,�V^/�=��%'t��K��`��!C;k��1��T�ݳx�bޮĐ������g���������I����N����Җ��B-���-٬5a7��?WϿ������[$�H��y+=��>4UL*3�[�V��Ͼ����f\+���WX��</(�Xb���	>45R.�-'-/��7�&x�Ԡ�x_��#*/e`�1�\o`���]ά�_K��uqxQZe�&�������S$�f:�֊v{/���#��ʗ�A>�)�"���jŋ��k�s!�B?oYa40z�J�3K���bQ
G �Z�db�c����D�7�Z�}K�X!�	����WAi�f����~����1u�A��t�lJwJ���[�^��z!�z2��F��;q��J}ͦ�-�JV&�����_l�|̀�^��x�P�:�/i�U��Z!�j2��O7?�*$	�-��d��/�抓8�:ԋ	-*������æ���B{=<�Z��rWM�}Y��q�[
& ca�����u��~�c\+Lf�8vb��~_�f����nW�{� xG4%�ٜT`e��/�����,(�7�����@�z8�����yt�r~봹C���o5c
�͝TvmiNM�?�@4����-}{�U+�~7n��%+W�`F���i
G�\h� ���_��B����䟥���=���F}Ez�H﮾���]��d�j�d:���1Y�I���h����ʬ��+���/�\�l5��؝�k�o��knk�Y�O��&���C����{mk����x���r�hn��vQ��Q��������Ğ�A͆����!J�:��%=%�_ȌjZ�%Z�>��hQ��u�����Z�x��:P�����T������J���6���I4�Y�ae��7��7���"�����ԭ�5�:
4y��hWf*���z/�����s.P�˅u�$�DK}����%2Z%�aB���8H�\���M��EɽP�e�4�Ӝ.����[�;�\������]��6$g���X�)�U�S����?J}�9���[����G��֜�h���9]+�ټf�f+��=R��~����[��.J��t�(�΂�]����vL3֛x7K�td��ʨV�Hs����ʧ-��\�<1�v�߲�|�ꂯx�g���*�|�IG��J�;^� ��uP#�K�]�쮔6�;W�F�u�uIE/tz���~�hjhm�u;,�xI*�n���L�|Ht3MC��'ԝ�bb]���)Y'��ģ��Y?��;t�R�I���]�^�
�{�G+ŧum�޿`k2���U��6�_Oߙ�K�I�c���2v��EaJ,���|�8�6�|�+]��+�<zQ�����'"	4/�M�C3+S�O�+�d>Wv��@'q)F��p�l�$jQ|��%��x���;�n�Y��VϨT[��KO�>�+�\1�5co�����>�Z�A;-D]���\�9�&)��5�lP�5̼0���6�&`L~6b���M�Y�ڷ��o�Ǭ��*�����a �ڥ/��F�?.�sm
/
�"PK��ӐeC�N����P�XD>J)�� �HVv(�9x�k��B���[�w�=��ȏ�Z���B5�W^dF��8�����S���~[RekS�yЭ�tL"�-zX{�4{;��,����t�[�pX���Ո�1G�h�:{�o���<I��2��{+z��9J�G�ǼZ>���M�jw�
���O��	�d�ɴر��B%�.�v��:u�\���4��m���w��G���Y�:�?n���_f^�7�MGU����W(�댻�����^1���J�������~LN{:��E���g�� Pnt/ⳇ�`�u�>���[�e��^���ֽ{�V�����������F�QYHȆ����K�T��yC�Q�[hQ'�)�{��)�x�h���{S��T@�R�q�[yB�J�����J��D��4�W/N���k�Vӳ>꾚�)S������:����PKTJ�����Gۡ�Q�n*�;$�+��Oqt�W���:���V��+�j�9n�OLm�������!b���Z+=@�Sl���D �ќ�_O�r�`�b�����3�{l
L���v��E�j����Kȕi����I+��Ϟ��v5���wI\֚��Q�+ӽ`���6�zG���F�㳫����H�3ϋ��G�h�=��G޽�c�7�E�P*<H�A���6�/�;����՗ȝ9���fg����
Pg���&�65���6�t9��y��W}~�?�� ~�{��`�4?�y_
E���4J������Џ�/���Pgs�-��O϶�d��E�s�s,+�u�Ie�����~cR�N�1��!yx�1�a>�?v��>�CR��D_�=!xQfd�oG�2���2���Z�A�������c�D�櫚�]Wq�	��xSI�k.�c��)����b6�v%?#
f�7�#�2e�k`n�/�5��2�_KG��";P�)�עB<X)r5�,��9ʘ�_�,^�Ę�#Mi�G�r�����:���}E?�1��G��%:�c]Yo]��5S�89Mb@ܬ�?S.���_d�^�����b���P���9/����uТyJ��0�8�h0f���F@����n+,�NQ��cT����?	_l1~4��Aρ&۞��gI��p��c�16wi���n���\��#���5VX��9{�d����-�P�,�]]^�$�T�T�`z��Ov�CD ��3�՜t�\����] ����5�E�t��ѿ�<�S��*��ʿ�a��A��y�'���5k(5הvuTй]$J�V$�j�{Ǽ�n�hnHԘ{�p�]S�)f���elq���_f��w�hk9���1��6Q�����gM�E�8�m���an����b����w�Jnהܖl=�����Dk.d6�;7�M��V��-c"�2ܺ4�v>=C��m���B/�6������u��mّ���s��LS�T��㱊�p����G!��B�����E�HeI�'.s!Y��߹��&?	�愈�+w��%_o��ů��b�/�Ɂ��GY����5f2o���L�9�M�a7��,��w�F�W�ȏ����:�ws��>g���Oyʢ⳼�&�o�����VU��ֲy6�s�_']r�[L��.l&ˌN��]�y�͡��p��	в2\�e�������O^�܅d[n���.��XI�J�>�noP�W:�F���8v�0eT8Z�L��&�|��f��Q�w}���?�\�Յ"#������:���<㿘���5`�_�V$Q��a}��N~�x�u���%0!�5��ȳ�;n^�d��GH.��?R�&�w'�1��^��U;�يDWP�&3Q�~'����,��O�I�R����J�ճϥ����>�ndxu;26e��)]l'3�q�������*��a ����X�s�\���l�U����i��\�>y}�Q�u�[<}�)[r!Z���2�gv���Ꮎ{�CKp̩a����g���-��Z�X/�Q��ǵ�_�&n��6.8d=)g�p��/F���9�8��b������|��,!|M���)hY�����x��<�u�	��z���gA�X��R|/�Bwd/�$׮p(b��{��㋥N��lY<��ao��N��{-���;��v��q�D��x�f��"{x��-���qՃOvz殺��p�1PD�}��g��ʣ�lo\�����]����8��TD����]��'�J_���H��H��Ϧ�Zs�����-�+XF�+C�e��{��̥<6��=���o/�����%��t �����	�#���OU~���@EA�*3�J�ǃ(&���rK=I�K�'msGGW��|����O��p�K�<�n �^&q��c.�8DN��|�r�o����R��pq��x�>:p��N|��H��t\�>�����i#�?��x�"��n ��!J:���˺^�N?�P�2:������1L]�(�q[��Ӗ�o�\���ϡ?d��e:t�%"��2#�f�U�|_7�?Yu�5r�c�����H��9vKr���^��AYxV�0]@��NM-w�^��nUݴ�f��YW��'���q�����+st��p�����{4sn�к�&A]q�J�<�R�B���ZC5���^����M�;Iנ�Y��Ĳ�O��7�5B���r̠���b����� � ���fg�J5q���Q���Ox�,h�� ��jq�%��;Ʀ�$^�8�1\�C�h<����_���f�bJ�6)������g�X[M�l|:t^��v~��w��%'ǹ�2:<�N�q��֯�&_�}Ǹ�_��b/�\��җE_+��6m���?Q�_�[��2P3{�J#<�o��m���5���W3��I^�#}��p�i&K�U�㏶�����s�$����5CG���*�l��r�a;��*�� Ԑ�:�)w��S�&:٠��!�g��lH�^w��m�rF�v�Pٟ���!}�H��*�S�8F�=����˿�9�Y&�:"�^�����{��p��p͵��:�I����7X]?�
G�Yu�Z��$ߔm&�Q��A*q��A�t��4�g�K�k�ی�S��-d0(j�+����//�T��J�F�nR h�(����&�@ި��Mb>#T{o�2K��6�1~�w22s��K���2 ���_��})p��ŭ+��&{�ĪݍWm�Z�,'�a*FC��F�����蛕m��t?���F���v���x������-wǅ]W��hu�u?��.�����G.c>��mC�`��|����D�bǌ��ZZ���<q�|���<�B����O��WH�d��Y�HA��2e풊0Q�j튷w4e�l@��շ�#�+u�k�z[����tkSP�	4g0v�o3ߩ8����M�=�Op�~D�
�ct�)��1�ISOG�8l�ՂS��i5A"_\���@�Jo�2��( u��}�~P���M���g"'���&���OƢ!U)�ChWԾ�}��owq�ߏ����?$
B����A[�!_�؎:�c�J�����$u��������y
'q\4lw&z��bR}/^��E���2�馅�Э����O{!l�<c�����Rs����1�����f���9#GU�)������{c#|�g�"w: �|���m������zL[G�KI<��:F)�3���?2Tc�T��Y�f^��x\��$|k��Ỗ�>I �p2
|�v��	cg�cy�sP��;q�;��~S�o,E����a��NN>DL�"t��W�x��*܈�q�~t|�m�6�����.�A\6�M�6���.��ŇD���������%;���YHn\��Ҁ�,ϑݝ!�� �Pi�$���ѽa#�zL��YvÇk���-���0���~A��>i�-S�V���jP��ȓG�c$a#[���1)�5�گ�?i���.-e�~;n[1?M�����ƌ�0�Å��{�wFg����H�x� ]�X�>f&TW�UjSm`ypT�?zͲ�oӶ�J�7��K��Cou������y��3wT���'�&G��Vq���𴟮.2��V��x�����$���W3�w�4�@L<W�b;��~�mD���DJ����]!I����`��|�M�F}�����,�����ʠŢ�[�Ю,�̀'J<A�|��%
��I��'hǉ���W��D:|`ǵ�+v���|�_��/*N��5�'�	�?|�K-��?���{{h ���D4y��������9�y�Q�걀��=�X�M.'G��j���#��4K���|L����p�rxr����145-� ��V�;��JV7���%�|�"&~zե��d���]���>��?h5��A����J����Q_�нD�*��.���^�H�B����W�ߩ[�M����\8y�l��uT�5��6�H�I،���0M�ci�7|�x\u�YO�N,&mR�0��m��U~��
��E�)S��zU'�����E.><�y����>���x.��w0X\�f��:`\lY㇩o�흓��h��O�	�բ�7��G�����qc�E���@aܯ1��!ݼ��������ezh��-#J~��l��mRKL*>��Z�ڦ�4c6�%�<�8s�H��*
%j9�''��*��(�Wsbb�X9|P�i�ҚX��wb+N�z|2��ʕj�ڤI:v2��73�0]����q�s!�Wz�yU�8�K"�S��uVz���|�c�E�R�
j�4y\|�cG�[յ���P�����BGR�p��� 3fp�d�t&u��,�;c�@[J\��,<q��ۍx��]�|�]�{�λM�����
 r+7fR=���
��I��������v�'�}�p��=����)�I��}�S�����&�D-UM�ӪvڲZdR��Ω��H׻��u�A����'�"����̑��t+��e����P�lΩw@����v/�.�����ֿq	JV})�
�4�r�
ް���LR.Y/T���M�-I[{�e̺W�my뭞1��)_�*�>����a�����\��4ڲ��G�llq�|R>���<��O ��M��d%-`���k�o���ިD�/��������E��p��s� $S��T{���+��!e��,�콡��oD�|������Gl���+v�}�y���)yw|�y�W���r
�zK6��;P��7�j��3�(zhD�E���r,���y���qc�i�*&f�!�C�r�p���.�?k�U��;کQ �����pp� �xo�;�=ض0�]�w����9�� @���;Ӎ��7�M�T���Y�n��r#{���˥���N�<���:利��Mۑ�̱�P���e��oR<#�տ���;ڶn�䯷�S�r�h=G��7�L�k҅��ި!3���	T�c%O%.U<MXIO�h�7&d��x��h����6�*es�%&q`��H�<:���!�f3A;ejF�^՟�<����a��Qg%��T�kUȬ.d�mS���d��l .ž��!�+ĵ@�B��҇$����o޳�2��J���0DF��R=�a^z��a���v��.#��������6���q�{FK}�����aLiNM�p���Y���n���+�gAA�����B�ܞվC�ո�m���p�⺫�G3���2��?g�<V�ғR���[��!;��xE��q�T�Kt�ם���7ji˪����3�Ucm�����B_��:g\=�S�������)�z8�i�I�;O�v:��˂lc�צ~"%`X1Z[���>j�[�a�X���]��|c�{�ޯy�iO��������0U����n����Ķ�	��v��Z�s�_���jx�]l?��KB�m^q�7u�p��Q��L�VZ'HW��}�0� >ݿƉP�����r�l��2�2`��O��g[6,�������i�Z�~�s��-�ga�\���x0y�Cts��/	�/1�]o��)x�ϝ'?i��` �������mn�	M>=_�3e�v����)���jۧU[H�����������6��w�U��-^&V��B��Q�m���q��S�7�x��^��;��Zx{�� �h�y\���čGR�.�%U��X^<��k�^��wX��t�M��ȳ�t�a讅��<���b7\׈�]�r�t-wo*���J�nV�Ǧ����%�V"*�Us⧣iX:rF��1T��ָ����rZq�Wg�Б  ��2{���7)��:��hat��zݣf�d���{�~:�8CJ6��1�>�=�����-� :	���g���AB�q��K�Ҵ0`�8[�W��IDJ��d=��a������	��\��r�D���J.���v���i�������3ri����g$C�R]>��ε�K?L��_B��,���.�#�aa�6U[Q"Zڣ�B����@⵵���sL1"��v�U������
u�L�������~0~OJj�e3'�j#\���7��!�'C�u��t�H���{?��τ�-�_2a��H�|��j���t����+SAm���g�������L��B�?��
�]'���HsK������z�۸ꆆt���{�C�C΃���ĄUYY)�qI:=���Ͳ���/�)�O2��
�_��+���?�
/��������쬠������+�z$�R\J������~�f�J&N�&��?��L����ה������<񎋋{����ϟ?�K�Q������o��_��צMFJ��Ƿ��54�588���������������I���ӭ���Y����< D�P_600P@Mmr�hݵT���W1Zfcaَ�Zw��۳}_fI�T�����t���W
�	��%%젢�gdЉ��A/���q��_d������d�s��`//���Fa/8xy_b��+!�韮�����CU�1M��6��~Pp����V,��蘒���ؙ�h�qy>GI.�oMk5�H����*�������tu��u%�u���3ps�|�z������y���̧��J�iii=�)��%��]�U�m1}����11$,,,o��dee������ζ�x;�'&T�ܽ+hbb���n��۴+����67���h����8�2�����BBB��RR�_�^�AG����#�����QZ/'��䥥��������5���NKK�i4g���srr����G�к,�UޠaOO����20b�Ѐ,���Ǡ)�Hll,����l�	��EES�kkt\�ƣe���߆��RRR���yx�PQQ��FJ�v!�Z[��)ıa���v��RC��㨵�,�Y¬�#@kA---Mư�'�����yxx�vV���K���=Ʉ�cXJZ��ׯ_�����{�!/���!;v��=���S��i�t�I�lXX =��Z�ÝU��	ٙY��4}�.����ڭ���k�<���1|1�;�?RR�{���\Y���n+���65�:<<\}u���	Z��Ey�O@�v������2k�N'L�90���ۻ�ׯ{ E�������_}}��������A���(�2���u_�nD�VP-�Uxll�#���BV�?*ŕh�v1��@�pNo H��Ϸ�l}oӎ��e��T���HK�#p�]3a��#yX9���W��QIe��\]]s��J�42��ۣ��e�@��:�@����^�@=���>h����N��U��!!�
ڐ��!��!�l���E�,����o���	�?�3����T�56����{HB�����n��iim_Y1���OD��{�g�HYEZ_Ldfa���Y.�/++��ۘ6;@�Q���+�3V�oml�C!~ [r�B����|H��A��H�.��2������ /C!��5,,,0�"�󑭥��@� �)-�FK�ή����:�u�+,d����}������������Tj�d��JK9��G����n߆F��j	.��P'�s�v>X|HD$a��Y%0;?�8�^�OL�XZ^&h"�q,��^�t�y�r��kbb�|qv+
�Ȗ��l���`���>��� <6�qŕ�s��ǿ\��gDD �PAA���E>���x���E��$vƪ�틽 '��ň����q����!111��<
`��h@8 �)q��w�����yX%(�����S9`>DT֫C8DDDf3�~��%�\�_��ZY�h���x���V1].�#��nկ���l��������5Q���7"�4շ�zE:�n5ut�������B*W��N����--��L��6Pd����L��FA�$ �
�.�Ä\�t�����֬�zto�ژSF��Y��cqY�|�M�� ���nܸ1o��=3����A�PL���c\�3x��|G�or�3g��\Xht4���WM�u�!��~��^A8�l��
�t��ƈEǭѿ\b��Sd4���z �08���r���Bө���˘t�4��y󦠨��:|�nZY���-&�Z�@gg=���Elq G�4
�Aap)(��:R+�d>�<���Xe[i���&�Tl�}gu�=�� 1�nSMT1^����Q�����ά���~�Fo�Ӊ���X-�yT�[�����Mf9�uk�T�ah�AA!I(W
t��\�~����2�ؖ�!0�Fo�,�W%�+��lE&��B>��;;֙$�_j��Z4s���JN���/r�&M���Q2�d98<��"vK���5]�8%���h�����b�ń  )�UN:�";�����"R��$�����B�Ķ�l��o��l�5�v�OH]S�|Q�o�xB�ݸd�kJz��=ZEpc�j�0�����?���g����@$vhHRR�s�~dB��挗�倨^?���p���\��j;��i	{�Hv3Rt"Nl0��6*oX#�W������f��xnf	� �")��Ҕ;U�����%.e�F�x�J��,�rR(��C �@����{P�82B����$�AzȐ?|�TT�P�E��G <�!#$d7��s�9��.g��4��c�� X�sA���6�92B�˽)��
�"��|��?AWf��}�J3�1;�cd�ƀ�oCO�ۮ����K^W�
�/�W�@b7����#V�ǉ�$#�}��l�+@����S+P"8�l|�\	� 33�⇻�YYY�Q�=�bttcQ����7zT�i�v��κo���ϔ�$Ν1ӗ]L����l�<���jH�m��s���Ў$IDLA�|SSS	�����@ ��J.b�t>Z���'����@�b>�q��l!�.D�i����]�S�B$���D������*do��������{�g���K�߉m졋E" ��^�����.�a��}�X!-PMVN��H� Y(x�?��x�q�-�l�0qJw��%٦�rA\�_�Ft.<7�o�䪀J*Z����nj�@�ؔzG4hB�Q��@��ç}���x�߶��C��+�V� ��I�����x�?%�}J�۹.�'��^6�' *�*�e)���h	/@<W:��A���I��K�Ni
�r�B�d�Z����f����B��t��E+q�����%�u��*ޱ��������zw,�3Wn�ȇB�-&E�ƵH�]�y���bD��:�GXX�%4� ��W��@�DbC ��0�=�N�~/  @DJ��?#�����{O�qŏ���D=}}pT�{��H]2@k/��'�#�A[�5P������7��A`6o��O̿��?i:���RYB��oee5b7A29��c%�@H��\ۨ�;���.�
ظ�Ȧ �qK�����Gj\�Z���!Q�c�q��|G����eJO��>%�������r�U�Oۉ�7�@�%"5��^넧�<�Ӕ�?p����Y�BSj3q�/!z��,��722 f�>�8�5`w�]�=^>�9+oee"ƐI9j/�d�q�4�f}�*تjץ�,���"�DW�|R��J��������7��{g��7�R;4�UQ�O�+ǋI�
Λk��Jh��f���%�\�Դ�I��O����Q("�'�Rח�%!�S}����\��{҉�W�.W�~;*1�ˉ�b�s%��d=*>>�ǔa|.U�h_�?:�755���5Ά����>2�?vV,�zo7tT~�}�엪!��V�1O��~^���.�Ls0O+�|VԌP��&usz� 5-m �."�����u q�$@���A����4L. p߽�dɞc�{��#�:!�	ӌ1������OT=��?$��`�?"ff��}z�u��Ua�e�PJޫ��f�+/Z �F�Y�
� �zB*����X�u��펂*<�����$�������ԏ�bN���;b�5<����g�RXs�~�-!e��(����'''��2�UX��&6�AL'g"4r����>c� �kl,�:���4��A���^E[KG�c��X����P���R��~����K�+8v2���kn!i��Y���2�?n3�q�{q�{q�g��{�IQ���d;���8�*_��`���TV�iR�P��(r�Yx�"��7�Hʨ$��Ր�����:*a�y�{wFx�������v���^y��f����< �H����7�*출��Q������ޘ>_�t) �Hӵ��NN��й�t����0������H/_�g��&rvP'&�;Y�`��&l����Xd��8�����`�` ������d�+IIY��&`�SҨ�n�&���r��IS���k�V�1KG��hV�l�+�9��M���,t�q�����:��8���Ef��������ꪓ���D"�30���GԛSCF������!:\���'��9}Osb�\�����@�ܗ9��_�sO�{1@6��$�p.���=?%�Ӻ�[�RR���+a�0v�5\?��ݟ.Χǻ���]��־����A6��@�Q	Z��FЖP}������Jx�<ռ��\P�������c�m���`�.��������+ww�m�ݶ�v�[0R�M7�=�|����11.�pZ��4��q�&<���p&H^��������l�C���1D�8������o����AÁ����j������QRR�MR5���9d2h'~{OKJ����ȷ��۷�Н V�Ag�FC�6f��l�_(�d���u�=w�0��d��h��f��o�'��߂m�b8��v%��bc;�?�������l��縒�o\���xy�_��ۃ�t��������&g�//.�1��<L������;-\�2h�~C�P!o��in_�=L^R�д�t
���k��C��P-��S��Kq5Ȑ�	WTVg��d~�ǠR�d�����؆|q:;��:є���}�`�5�)��k��#~4�>}����퍍���l�QX��p�I�ËA
ak]��ޯw	�nvo��ת�Df�E}ct�l���9R�sZ��XvKl�2u����Mp��I��xZ2�jWP6(�m1�n��t�rw����h/i��7�)�������o�6yBOS7�+�,������TT�!�˪��!L�U�lnm�T��T�d��������׊�HI%H�,���<��( p�;nǯ���8�J�=9�^�=�'=*`�a����Vb�Je��ὸ�#>�A!�܁qh؀-1 �����f,H��h<=<N�DNTA����HquRJ����;��v㛱Ľ��w8�Z�eV�!!ɀ��n�� bCU7i���q����hI��Օ~�W��=t OQ�W�	�V�����cqQ�3��~ Yє&��e8υ� ���:zqee$,(h���������xu�������&�.Q�_�vy�� gV��t՝�0�����ifE�0@�_�����;�L�W��<?i�>�Lp�bu$I�ˢ�9����;��o����́(t�B��`jT@�Ò�0��ls��ՁSY��"� �f�u:�V�
�W��w�|	�������C�t������恶�Ʒ}	WWW�6�-L��
�S�Ӈ v�m|�_�,^s�$�X���xy�!,������PP�4��hֵIsS�oHʣ�|�Y���-(¸L*�z��M�Rʆcvy���p�䒯�r �����Nz�{�n�D'�f�6Yi��i��R��[dÙ-��gp��>�/\���1��;��c�1\��y,jb�>l�F�y��nk��5i�g�v��j��f�u����N�P��Y~��U�Г��N�<̉ezg����Ymllܬ�F�K�1����Pu�Y�u�ǂ��y]�r���&(�������_� ͏����O��I7K�<���G��N��H	�$,8R4���h�ٴw%}|�y��3��b������q��[I�2��P��4Y*!D��k�2kc�ne�HDbH��%c+ً��3�g�>_���3���׽1�<�sy<�s^�3�w~D�4��h�ĭz}M�x�2�����4�8f���w���8��3a���m�H�F��t�_����xtz(JK�͍H�P��e�ίc�`�?�w �,��'�̘T�\I+�Ǳ�w�Z�N���>��m�R�`^�4k�hR�Vi�R4��"�4�6�[�B�RHܞDD�=�kRXmS�Y�������8����d5�/�u�%�Ƕ}7�_�\�$��>�ӽ8�|e4�\S#j�R�A��)�� ��6]s1Zk�֪��^y����&&eQ�\<O�H{��F�R_ig��Nt���Q�w�H�-@^*��OZjϐG13U��˔���4"_"����τ�M�G�s9�J��R���:s���M�D��r����=87��\���g��������pj���r8]�5�=��=�3g���IV*�F筥T�\m�SD ̮A�����T<���\�[�=�*
~���1�V}��D%Y��g�
獩(��lCb��H�~��2S�H��Щ�����]�����)
Y�Vtз��e~���B�$� +�7��w�r�[�|���?�̷�	�.��F�2� �3+Ay&&&��q�*W�F"�uv��ފ�e�D_H�,IE��^�����\���'�\��k�O���N}`omkK�Gz���a���9�X��ˆes�ː];k�{Y�0�w�'�ϸ�~��*�L�nQSW�^u�lŀ�;�+�����%���>�8����y�E<���O���=�Z�m��NM�T0jeśM��4�*���a����H���x'�>��f��BU��B�1��4W�����o/oc��g��
]F�Y��4^�J�o�l�������g'7z�TKSp����O�\cD�mj+}�'����)c��q�J;���CƆ�0h�c��!����L$R�.R@�|}i<7�_^�C�N�M�H���n{WL/��@�d���s��f[��FN�CG6عkW���kFJ�K�l.`���_}f���~�W���ȼ��0��uH�/�qp�$SO׷��)�}(�w���z�
?�}��#M�fb��<�g��`�2jaϚ�}2DY�d��1I����s�o�&�K=�T�7&���`]�<��S����� �.��@�z(���U�<4���F�71C��鈴O��� i�?�������o�6��'���<��s a�6�k���A�e��D9C��{6�T�c�#���Z#:�`�onv��SO
������L�|	�y���(^a��v����1��������(
U��
���*QΫ�5�Y�Dk��F1���<����;���5<;�F�7k�R�eJ~��* vuuU���=��i��i�������UK��J1v2���cTMM����ЇE#�)��*���%�� �ԩ/�L�˛
P	��t����6a���p;7O��533�rqz���~�f��k2�|#�J����ޞ������5�pQ0�"��{�9�G>N��l@��1��V��??�J�;�Nմ��">��׶�$�;�{6�o���kvo��G	E}k7 �@ΰn��hr:�.y����vi�P99��Q���-rqȞ�8���|�����o̽B ����:�rKF�����>�&��s�A�7�.!n|��N�Q\g3+]� )A���� lP3k� Y��$��Ԣ�.ʂօ��lq|(�`�4ȸ�J��p��:ُ!۩�Nmmm�>��_�e�n��P�~l���g#(Q�O�>�k
��eo!T��*��z���(��G/^�S��\��i�q�*��<e�R56�d\�o}E�6QSS�kM#sn��|��5�t�$V3I��<�%�Gzz�
���w��V&������ˁ���G���I����F���Ȝ�c�N}D�>�  Ѥ0�P�!+j��5ccљ�殦�Ǚh�6��b)����0'��'�so�
����/�]Ϟ=+����և�!��%j���F1�e�;��!Z8߲��6E�C1�m��C� �����̑��h�r�#_\��xV]�*��jm���E�j���S���u��Y�H�W�5�秉������X]0a�P����8<4T\��7u�f*۶��Q�l��՚�A�"G=����Y�������(�I����OB2�q|�k�7m��45�=#Z����ː�x ��vv;K���_% j\�P'=��tܸ�:=*�<^�dّyc쌼}a�X��טV�-�l;�rY��]����s�t��'�O��ݼ�m�j�d�왟�fU��A+v˵ �h���O���b�a?~��I[����.�x��D��⳶�������ަz�.4|��0�B�|���v
��0,���X#����&���f���p�ib1��B=`V�P�_-)*�?�>�+��2������a�w8��	�g}hf��۫��m��O�2I���sJ�����QBZ�M?��h/���rJ~�E[�κ�4��������'�m>�^v}�kԛ^^u��隚:�yz�H�IeK,����ok�Q��`Ȣ���Z9��_���>�H� :�M-�B�WV������W�DЮ�8�Kt�X��G��/��5�>h�Ħ��$�oBK���(���N�|������BX���DWwa��tB{�e�CC����Os�^�O�� ($��'�!��o��O�U�����{Ё`蟷�%(e�����r�6���S��{��%�3#����5a��ZJ���v�!f���1T�PU�U�u]�Əq��F�(1���x���.^vm�qvaA( 8�7��OMW2�酟��0���3�9VWW�ἜsW�z��{�Jۻ�����Y� fEc�c��j�ܫ",$��-\��FK�tuq( \
t���A�%s��/<�rT�<�����z@�j���V�lcmpo�O�>>�7�|�|Ｌ���v��ɽO�r�榦k|�����:9�uwq�y�}����/PTB}���^ qOV`ۖ� ���	�����퍌G&3Fo{z T��X_����漕U��s�a2gNu��>��l:�P������<h�uC�Omv��m�ܜ�X���ma���1��y��/jX���R0_qL�(�t
�!��ý��au���X�1.�:s����vq�����h#n�˔��bc8Z~T�j�+�x��-���y�`�	% <�I|�O=G�1���	���2�#5�t�f�m�3��W�@IG�d�+��~�W��"�<�Z�e/K��S�|��. ����*,.��D����K�姌��)MrB̇��d�q`��ƴ<;e��㳓��;�*S/EY���2gJ'T���,,gȢ���S� ]H������#��{6M��1:6VHaKjW��;(m��JQ�����7�� ��@���被n�ɳD�&�H~^����u�p��e-["����|P�S��Ah��t��Y�q�B��
\��Ŭ>���,w�������<]?�/	���8fD�Ѿ|�!�k�����w���O����O~�����hoWur�O�$�o5'������#˫KKK��C��>*J�G����<E��h���@W��/��h#��^:�<�9y��{?��^ڸ��R	B�s(��L8�e����x��~q����\74\���6��b����yR��"19��ܵ-�N0Ѫ;n�z�m���*Y�.2��������S���|1��%�����	";�y���y[�J_����{�,N �~�.���3?&�����ud�x��s4ٰ � nkg�D��o4�ܠ�xf�4�W �]�i�o �t�Y��`(��`o]�ZT4�vW�^;�$��:tC%��V��EE��([ܯB6�#̔+D��,*����j#_�f*�^����_cS��S�;"��[�@%��_��ŸFU��6���3�$$`������H�v�f��5pc�����g��
E�h+O<����Pm�4�H�7F[�`ᴐ' g����Ϧ��+J��İ�R��T�:��~ƅC�`z�U���9��|� �C���g?�"˵u�z]ʁ��H@��)a3k�� 9y��g	�\��uc���H��W-䷉��'h���y1�DU,��a�?��m?5<23'g~V���]gOլ\����Q,y����|��V��Ͽb<����Ν;� n�.r��Ç{l���ss.��	)��;�O%݂�=nR�N+7��%�����@Z��$���Lz%�򎓝k���c��S�~d��&�PX���]��fy��#��h��;�����O2<�+rL��j�=����kܶG9ܵ�Ԍ4,�O��Rn4#*�~�^���
���D�ieS�����܅`�n��5���Yߛ�7�7Ҕ��;��^�����_�d��O�<R�?�R	�P�}c�&ƅP=H:�A:P4R��v���т��J�1&��]�%M��jb"��E�K#\��c<>/�v	C����k&���BC��?-�,g���rbGm���c�w���v\\���=��v�<#C$��-��U��y<�;��ˊ�����m�>77��qc��߷s5*x���
aF��,Ot�X�:1�x�:R刬��
ޭ����_dѪ����q�e����׎#�ra��eD��U1���qy�l*E����Xk��L�ɫ׮���[�x<��Q��l��֯UA�I6�ϛ��ǘ���w��#���,��㾇�i���
"�������%�"�Ǹc'l��JI��2��n��q�BU�V�Y%�E�7]d޸ߙ�����Y�N�b�	�/_��d:PDH��u���e�����@���w~���� ^�G�l���E���ۜcn�P ߄~h��2�
g���NX��H�%���M��rU��s,-�T&�"�C&�?�lQ�lN������_���m�!EX��Y��rb��rK�E��k�V�����=J��)n��e�1Kii��89�B\͛��&�������o�v!��sc�J�5���M�\�ĭ�ׇ�^5,<������DWi���S5\�X��w���.�}I͆��111nn_�2`�~�}O�MI-<!+3�1��鴐� �O�2j��%-�f]� �ʩ�f��D�Dʛ7W�/�m����
�V���|�*��`��<k��ړ�и	sp�xG�-�x�%�5�V���WG#��J�����0
��K>��7��i�ܘ{/"����ҁã-){&�ʖ3`_bCC�:1%%E�dq�3Xݖ�y���P�׌���F���m�����k��'����=<�7��a|E^SJ��3�I���2����~�WKu��ڬ��wbI�B��vz��+���`%�`~����d�]��8ت.ޡ���TpL�uI�v�5,Z3<T5���{`P�!s��JS��o2E�{f����?�������K�z��4����k�N�e��",�%��~��2�`��7���V$1*�A�������_��Nbb���ai�{d,ha��p�G� �q���kVa�3��%�a�Ex�P��|MQ�������S:P o�I7,/�+i��&K�Ƒ5�f���_�� �m&md�Y��W�N �J��X�N��l�v�����@�,p�$�VVV׮]{A��ຉ�Փk��*�����[+"ҭ� (�
��ajf����r��ګ�إ@�ځ��T*������d?r� ��Nt�[U��"����C>C\��L��Y_=�ptQݗ�eЪ�[�
���:��l��[��<I�-4������,�:�;a�W�x���x';2A:d���09�	PT!k����T]��&��$� �?�<:���7�8�ک���6?��2�#���ES�/����5�k#e��];w�� ӑS�h����Wd�����<��u��:�yt+??����j�����t6b�5�� %�$0���x!�a�O"~��k^Q��j�%ٺ1�������)� .��Ǐ���g����:��r�F�s��d ��E&%m<��iql��V���/Rn�ğ)�B��FZ�*�����'y�N�U����Pc'K�spT��.ZƂٷ>=K�K�Ka䡫
=��I����CV~�4�
:��E=꛵C�#�f���'s��Q��P���ty;�%�ԛ�6����� Rlͳ���un���P�یx<~vUO�hZZ}뫓����)�e��8��M7�}�|�E�S[�����	42�� ��򭦄W���6'�RZF��̓)0�9ҡ&gP�6��?;��I�=ʥ@�Ʌ�S������%e7 �1m�c�V2�����G2�� ���̝���2IH
����̈�T$���,|$��G�y��='����C�$�yT-+�8dE�UF�܄Q5A�ֶ��X�Z���	o��wfW���sP��g8n�CI�,�DyV�i;V����k7n��%�H���EB6�Y��̙�kE���������� 1z�/����Xc0�<[̼�����dJ���	���q�^��jb�hJ�[֧21:���ڃ[1��jVonc����M$��A#���$Q���mp����W�n F����n����=`�e7�|g�:ۂ�������y���x��Űz���s� 	5(�d��y.8q� Td�%�8�t���}�T��W��UTT ��eff6�ã��W���HÅ (G{z��� �}�i�L��ɕ+/^�H��v��~���	^�m� �Mo����[�����<��2
�kG�s�G��iy�� #Ҟ\��T|�F�2@���S�13�Z�VZj�l9�����ya��|+��0^�n�I�y_&Y]\\��я1���~=�G�b�(]]^pC�F����l���?�!�4UC$o�xjPZ������N�w��r 	����d�djNN���v� ����:w�X��ٟ����T���G��3�L�{��J�H��uXm��G���V&m�O����B�9zR��,���?�]������(#��]r��n�-�V�}��:�!~���fr:�,���`>��4����8)i2�Bu󘕆�o��Y��Gɻ\9-x;���#Qj�0V���ham{`{Gǝ���)(�OOOZ'D�C~'�]߷�٦Rq��O��e�p��0[Ȥ`T�K\���9�� /�p�j�W))����K8*y�V�(�t��5���5�����/o%����6l�[ ���ȏ�Թ�2H�_w�;�LM�G��.X[�T��0W�j��u�*�h��+�XYQtW��Uj`2����E����@��[�M��j��i����?R=w.�?�x�˩)�f����Ic�k�.��s8*LRy�$�m�ޫ�H�~��8#��߱���ׯ�+�����ǭ�q��5�������,�<�S��5#3�d��̞���!�޹S�N��'~�t3���Y��2�����uq��J�,#�s׶4���]:q�D�ZW�J���toy3Ԝ��ߠ���1�PZ͈EI��0"r��-?���L7�_<�������J��/�vP�d!@�q�D��"D��9���<g�����U��]�1Ӣ�?��5㮍|����zO ��A[��,tW��i~��?
��8F�{�}���ȸdm�t�I���
]2K���g�x���R�S�+[�к�d$���r`�0����{�E1�I{x=��b�E˫�]�.rJ�W��rB�hok{{�d~�d��(
�9:�^*2�<$znv��u�C�szQ���K��	(m��ã�h�� ��.n�S��_�t��khx����u�P��" �ko�B3i�O"�˼٣�2��R�H�Ѵɻ��`��v���|YZ\]*���<�ӷm�[~���0�vf��V�"���֠6��Q~%:�*)q�z� y��]��u��̼L�pe��z�X7'� /��E����#.G絠�P��'D����0I\S �4<?B�J�TRP�K�������F(��5^�tY�����|�m��/�_O�P�TR�0�ͼ/�������cq�HkE�Z���z/���T(�5��'�4�]���޿q���Ƿ0u�!ވu%��V�ʬ����"�D�S���q�K�J��]a���]~8ܼ��(22���w۶n�oj�lR�'����9�=��އ�y|Pt?mN,%A���V3nm6�ҧ���� [���O�Z'�2���j�r2.��lkk�joo�'p�G�E@W�6?"�y��Z�F%~�7 :��!�����ф��I"US�h��0�t�wX��T$It�	��s�Nt�dbb
�ˢ�L珁����8B��@�Ώ��H���EFFƊv,� ���Js�ː/Z5c��Y�
j32���.%*���#���_/E|�"
����*��33�3�nRG�|8N����V��Ĩ(�ߡ�ӛ�u����׊E��w5A���K�VI�{�:�|F��������rH��Y��D�L&$�C�rJ���;��X<^������� �_�5.�z��S<���Uh���y����ge�N_�.�}���d����JC f��8�VV����*�z�E��Z�f��[�?'dG����WRS�dr�?kֳe�H�э�t�B� ��C�E@�Vg
���l��^�"[D��-�#��#�7��
"+YOWIiIA\.��l�6�n^R�G ��"�{���S��Cm��a�ho$����Uc�=��j���d^'o'�'!J������Ĉw܅�r7�9A�D��Ob��7�S��b�r�`�!����߄�����*u�B�-X��<����[3��_�p$A�-���%���T����߿�wm�N4R�P��̽%�T:u�X!�Z(���4�}D|�0�����[��I�3���n���g����؜ȁ<"��&���������v��0�k�{�؛kt+���L�O%�-6 �n��v��MD�$��+�=2��\n�<�XeS(�(Z\\�Gy����)�$pӤڑ���/lI��&tD�"����7����tGv�/��!��-'��?��ӕr�.񗾾~o��0=&c��>ܔ�:l�8�N�8Jb��L��H���;;�3wU�t�p���,��L�q�c2��b�*'3�Tme�?��o�F*�����~b��|t���׬�	]��~����\]�}�zK�W�Nxj�ߣ�O#����e���������t�>�*�:���pi���į�`�j��w+�>�l�y���=_�-s�n	{��N�'���p�������=(�rIA�
��wT�v��K�<ʀu��P�e��ߌ�0�����Ţ���nAgG3+�!�R>���A��g�!J��Dhz|�����S7d�|��,�)+{.���G�*�+���u��9���L�g�X-�"H30�(}at��K|d�����9�M��{˥�:k�/8��2s�T|l�?��V����]��������8+]- P�4��*bӕ�5P���Twz�]S��X����a�s���"��G�����|H�2]�b<j��$sJ�u����
rV������_�
�i��������Gި���׸ty+���7f��C�ִ d�ݩTѽ�#5�S{��o���IX?��ԖJ
5�'L���O#�,�Mܿn�S1i;�ѭ]f�!Wݖ�>����7,�gr/��y���T4{����"��B7����D�rI�#i)V^Ia����Leӽ ��թb�	!|F�1IB>)b#ǚG�6_����g;~�|B��4y7�E�~L6��R�󱉒���Ns��ň
w��c���}��N���8��Na���b����.�_\	R�O�KDߦ��,p��Ɵ�lM@�Ո*0��EDD��H�6��6����8r��zP:""�|am��V�`�׎C�{��8�f��jok�{�����W뎃�{5)���!ؕ��Ʉ��b+r2F:���R�Vzt�ܼh���R�9�{e�dEy�`�ϭ�m���t�Z�����p��a�ӧ(ss�,@l��Lw9%%;}4k�+�9�Wi8� ���XsT5y75o	#�y�Y����}F��r<y�$"�冇�����_�b�M?0����-�k%����6Z�v��c�_&�	%��P�Ge?H�68(��ݱ�9���R�l���ދ%����⛶�M�.����]n�o0d����+���S]S��V�P۰��\�Z��8���vF:0�7Bm�Z�d9�U�VY��c6�\|܇Q�a��T�O����^�L�,��.F��S��z�q
vA�����].�,^iwo�ڥ毎?/�Q$��7�R�G���9��y���P�8�����[1��^I���۸�3��LKRR�w��f��fs���x���5�~��OcgD��3�r����۷�.xe��ҽ����hr���۷�>�����-��d�{��P�ڑi���x�b��9:b�i>׸o�ԕ�/}���h�v�{�e��wiS�Έ�w��e>;s�y }��@V�C�ܮq��M�B$�����9��K㓲�'��Z5mt7�Ȱ�D��p�]�'�{��e�v���A�Сsm�;hf� 5�(X"N��U^ /����C�ꃈ� :o��=rFH��w�5��^챍��$H�$���L��u��������'1� ��A�����
�l�l7�%�~i򓄄���e�e&�����O\��i����pllR���r������亽܈�N���}m��4:z���;vިʋߒ�_etc�#
I��$!Gl6�3/ڇ�M'�|\?z$���h��[�������9R���e5+�k�`i���!���_Z���4��S��8i&�ӟ ($D
�Ç�y�EOE5���ngMh�1�0��*�H�+��40�',A���k��7/K/�CF�իW7QʊH�~�����,��4k}��ݻ�NMCc������e{D��9R� n��c̛�N�#G��]�V��/(,,����s�M,����i�X4�lиGg����B���!UA�5v���Bcjj�:t�/w��y�(�Y_;d)�|c��޽����AHH���yO+�&��ą�KBZ�х�� ����b�Y}Nl#������8A�O��!��v+�V��zU?]���]���q�QQQ�PZ.+�����;�<�}Sa$)-ݶ���- *��+��02giɓzO,�(�<�����c5d�����Tf�SoU�>��^;�JII}��L_ ������kjv��:L�Y���z�{{�SC�=oĈy7Դ(]�4��)�`��ꊐ=�+K�0f�~+�bW�߾HF���GP���5��q`�)ZC�dΝ��ՠ��U�aE����E
D���> �����i~P�a�^9n7E��qT�2F�����%�G�86�V@lKj�A�:���w;V�����Q���j&�NƷf�ut����v� ����Q�ƌ�o}Dqpp��C��MǸ��@�9!#��&@gWWR(�r.>���fkM��b�y� ]"ȿ�P��?��oɉ��n��5���I.Q��y�e���7��
E�8&f~?2n4/�=F�5.,�]�8Ti�4�kj��������H��߻wo
�"��x������������ʪ���b�̢w����qjx���w��.NT�~N���tD��+1�����c���I)*����S��xl|��c�;͠��duy�;��kUP{���i*��-��W��~H &�\��H����'N�Rsqy��� �7��Z����B��4���^�t���F��0�[����ȏ��r��t |�'m������[O�"E���E*����(!-��\�n��+r�Y�!�|�.�SVV������w���m�,j	�g�qp�hA� �*��t����ƫB�`�Ksss� K�.`0������`c�/+ڑ#�V�����)	p�����'�j\d��X�KKϲF�"a|�t���Φ�G<&�
ZJ{z��I�N&�OCC�3�!{�����$��t���\$ާ+(�/��cs����g�!	$a�Q���22n	=�NM�X�g�؋��E`�
��כq��������PkcE!��<����b}t���!,A���k�ܹ3�'����	�S,�����'���<9��b��ǧN�jjj	8����a'�Y���{��in��E] ��-�L��:���#�-��"}��m��OZ}�W��VQjLJ����ϥ;����e�r�Kum�:p]HS�\�VE,���h��(��vgΛ�w t(������k���Y@
����H��!Kx-�:4G{$P+��3�,��ߟ� E�n+�H̯
ڣ�i�0a���DD*�����DB�"��~�����@&j��}���Qd��o޼y2,�Ғ,����/e�ŕJ�};����
�!)����dv4l�Q��>x��_a
����$eV�/��\��b���jԃ�Й��Z��tj�}
|�����zIU�Ȑ�E�?^�J�<8�OFVE��
0��{�וR�������y��%�7��{���e���K��%O�%F(�?9y�ٗ)Co+�WUޕ��&�tkC���/�jb�'. 0��@8A�f9)#���S�S�("0.�k�HKN>���M���n!((�+��߂���횶vF�5�8���Y ��{Q����4w�ǚx^J�]�����?�ܤ���o.�L�����2�`)$ pB����y)i������������N��r4��x5X
Z�٣ȫ(�T)��em..��c��6�>���O;>�u-�SّR��p�o���!ix;����ֶ�~ z�I(I�O,�!>�����WcD�@q���O��"ty�����g�n������U�[�˗�1b��g��Y��Б��Mr�֊{�1/^�O�p!��؊U\_����yd��c�������3�?�"�L)�s�������ove�[˂���g���R��s����GFG�>2G�9y��,��8�u6vv���aV�������fl��o�`	������_D�N������USq��C�bb1#�^����
.�z��`mc��|}-��4
&4>��$���̢Xĝ�<�� ��8�&�}hp�W{����U[;;;��V��B�Z�K����\�.S	m؀�"m���Oq5?�uZ��u��^ּ��4�k�F��*>�VA��GC\rqqዾ�<yO+d�r?�_�JQ��1t(�s\���*�,�W*�gϞ\~�(3��,s{��LW����9I\Lw�7nF�o)�t���_�PL�E�m**ߚ�|!���̋#����3��Yh 3�|�0 Flg�5�7�wre���DZN�f�n�t�B@I�̾�%~���5�;:�~{J�;w�w��λL�;O~,ZM����c�:{h�X��ė��� ���sʆ4��	@�R����8�<	��C�U-,RVF��2��JY�\%�.:;�_��iЭX�qICc_���M=.��g��`=|��CjzzÃ�"ŧ�{Q��}�'}���Z�����������	]ho7����o�m���hvm}m5!g�j��ٸ�z_n�q��/�!L���l�;uq�y����G8�\&�Ŷ���R��U��N�ɜ��x�?u�\9��X�5�n�Ժ�sQ���Z�L���U���ڭ�"��O�KN�,j��9������?��.I�z������6<�����9Y�`R�����O���64I���vmxc^VXX8	zh��L�Wg�H-�j2�-����!5�%���G�0�������d� 4���5�k���5��~o6��퐼�{�\�a�4C���NL�Q�5`cM�gy#>��h%���B�U�a憎�ܥ��;��3u���B�r.,�`��/vNc��*:���[�1����g�e�:�B�-��W#��La�l�փ�е��*e�K��X(�YD1�Y߻x}w��6�'Q4�p c�H��/�w�o��f�?��c��)��W��Xm<ӧx��4��]���mjI�B
���ĴN1���w�@C��4r�znPZZz8��w��ho$�Ы���P�b��C�/W�~+ME����毎����j�\�����t/��Ǚ�N��}e��C�_���LJNV�I��~�,��� �������u;j�<�t|ˡ��8�-��. ����i�_��y�jj>&9ď�2T�!8,|��Dk3r�̋/�vl�N��hD�9��x�ۻ�����OmB��e�r�tu�6�E�u?���xP ���wy$�.׹eWhj���>dNs�;�c����Nq���W�z��� o�>�����]����4X�֣`J��]���T��ϖ�֝����œ����.�_��̀3��u���h^�MJW�9�������_�.�� pw��𓗑w��WI�-746�&y7�O��9�O�C'ΫU��8�����fh|��6C�4�i���8N2�j�K��J����u+�{�߲�H�guh��ДC~�����ŚC.���qMO�
hU�_ޘ�)�]�3^���'��:cù�L ��&�h�c��+ĕ�F�pJ]E\Ԓk��S*RՒ��V^n�,E�4�K�����Y|�	fY�`��+W��o�" 
���JYfa���!���G�(<?��u�~[l�N9ԟ�n�xy����!j��&�"��MO?�]�W1C��[�$���>K�f/�����AJy[hߓ�w4	�!�K�h^Gq�� #��O5�����c	�:�G��s�[����xYzv�'"��7-,���\�`�H{��� t�����e�};m��ݸ��{Q���"���v��w{�RՀ��@��gfBzz�E;�h�*^��7�}e��4��#<^y��4d����V�Ϥ��X.� �������k�3J��Ϥl}nȝ|e�E�Y|nY|�0ڍ���'��{������������N��f�.#Me�@J��-�͑��W�k�r�^ig4�
6�4�U��d�C���F����%�ѓ ����%e�ͧ����Ҝ�E�'�����P!����.A��������`��ꢺ�I� ��"	�����������cp�g�l$��+R]@~Ǩ�4�D�����m�yOd]�����L���E�a��XlJ�<h�=)�m�,��y�y�<R@�0/Y�����G��6�rR��'��>���`�7�K����E��$t�H頍f--ynl-��_�Ԍn�m��|�ʹO(ɛ�@������U���+�G���Z��Q�h��/�s/����]��JJ��~�mcG��y乶}=��?_�S/S>�{#��ٶދ+((��k?�D��q�G���sR-^�BڮX{��Y�Ssaۂ0'�[�F�_�st�};��%�9��"
�j|n�@������iv�-����$5<����x����7{� ��q�F�r�:�=�x�V���j�V��zZ�]��c���]�H��J��"C��щ���8;�1AV�,�.F���7����!4��I�����e�#"�b��sd�
~zz��J�@8������
��&s��O�yN�P��}��ۛ�}������/�N��,�^S�y�r�����}�ۑ����I3�=��e(�P���O�۬�1W�˗�'�"4/8!�~D�/_���Vde�on�zRl
�dI� f�o�v��؉�V=���G29X��ZG ?`�@�k��.�y����l������E�$�:�����e*Ѫ����_��͆o��U���L��=�������� Vz}�N�ɦWf��	N|�h��N����ݓ���6�¡f�5���ڐ�`mD㻻۫��>�#��Mrs�sp�;$���^+o:kh|܏<w���BDH+��ɫ
�2��ow�s��'���222ttu�41$2$���a�1�K�m��\WJu��>y򤐏���sήx,=U�\�S���u�E-��
Y?��`��mpx�}���������r}�D�*�?}�d�9.7Y�^�=��u)��9�����!�D�k~�������5�q���g�5���H��<�P���I硺03�__ ?Nٌ�֫����?��x[:q_l�/�>��Y���n��gF�M###s(-��bO.�dQ���~uq�W��"x]W7h��T�A>��B,{q�ܹ �>9^"�@�C.b�s���h��r����o}�o���u�s4�bS��N�ss{�����-�哴GE$S�)[&
�!�dm>�F�!0�<ҀN�͛�U�`�s�&�bii�"����*L��c\`�x����j����8�����o����"}}}�3���2_�n�S[�93B,�]�ѷ<��2�_�����H����6� ���S�V�i�p?>y�_�T^����U�"���0N�@s$�?��{�0.Tt��y��Ok�z	�4 U�Tʖ�ɴ���S�:urs�����yJzl�k��C!�̾����9�q�2��Kc^g�
��ȋ��7���s�?�C�=VX��(�� ���/{��m��~��d�'��Ĩ�8ᴴ��+Gg�24⾵Ӷ�0O�||�}��-��)]�v������h2�1`�����F���Ah�|�X��}�wڪ��|��x6�>4����H�Ƽ����@��Y��E�cm�`xz2�}m�̹�ź���S�ϳ�/˯���@����a|΄pg����|ۘ7�ɓoJK��i��K�������0����s%����oIB��=<<�@Bu�G	YA�*�,͆��4]_��h��/�_�Ư��J :5?�@& טY�k7'z��
"���-G?'�9����V��l�L�%��\�04�\XV�,0����w�DXC�XI.�
T`C] �t���ڳ;�]�.�=]��Y
e�	ĒL�I�:)��)l��yG-�����q@��]�����pf����	>v������;/iiM��Ŏ,vi 
���-��+���e�b��/��[P���o���x����B�!b�]���0�Z�p��y���WIۃO��:��	h��O���۬o�Q��(Օ�|Y�}8bW������z�8��@��]�bif�'�xL�N���e;y	R�u�8�����.S�+P�$p�
,�]��A�yIC�(r�f}]�h�,���yL��iCV����AC�ӗ���r���;���i��Ou;�z�\�t��5'��dQ�h��鋃���*Ct��`^���Ni�p\߾{��k�0m�B�ޜ�i��E�\��7o~�����X<��\(�8�xQY~�ԏZ�H�t��3�~��!��r�s�~#����?����%���s�"�.]�Lm��Y�׸�w�a%"�v֗-�(�/6Wy� [1{�����Q����FfA�5?γ�}�6�����d
�Ү���/��Ƹ�ñ�U���A|�G���ɜ>5�|*ÉE��CCC̙99�_�=�s���"g��<ʝ�`K�u3o�i��Խ���Hq4�ˊ_��5������-�黺��U�b�!�v��X�,��i��_O�5׮��^��F���^�oyS��NB	�}��1w����Wo>�.U�o�
�8Sѯ`��[��������-DHSӨ6s�B-R�(D����>H�mSƸ1�܄^XqYKK��6�B��8�?RC��][|/�!�c�d��m�2�$��p��Ȁ��װ�7�~\?_pB�X�d��?�RΪ1F��6�(�F�o(���˺Sy^[\];κhebb�2����Ī-��F�/�c\����;P˅DQ>w�ߧY����_��;#�b	�tz��t��S�ۋ]���oɭ�'Rj�V]�+p������~$9���T�����HR,�*�G�3\d�+~}5G��7���vq���P"gHMK��nd�z$iQ\;8���;+���`�˗�q�.�]h��O%ɲh��w��P	G�ܚ��b��2H�H,ʇ�=42��|O��W1������;y	��L7N/��b��Z��~�����VQ	X��<���v�{�5}�. I�L�B�$�L�#*����7�$���8@�c����)�M@:�5�������|����mʝ���������T�b��a�j��J�-)���@��_�F��7�Y&F���v
���t�)��ĸ��r�)���WL-��- ���{�jy�.�ďX@��\�/~�`�R���f�,K |�[�E� ۟�>H�ծ�����m��$�`: ����X�ȒB��|��^�gϞY��0������jJ���\}T�������(������ҍ	�"�-��e��HJ����t�tw�tw�� ����u��z.�>��޿سgF;��:+�Z�y��~p�7�|i.��~�E��ƿ��qٕo��|r��J*nJ��Iq[;"�{��s�<���*��M������(�@H���D�_�\���	�dk�dv�^G�Z�\؋���:ת�j4F��vMۿ�Yt��K$�ŕ��h���6{�Ĵh�o^��4��1����x�y��&����Ծ�M����⼛�<��δ�+��]�*��7�IF�}.s��4�R�{N̛s� ����`w�+���2%*k��^�ay\�L��:`z&&��$k��8�ͱ����-�~�����{���$N�/_V��8$z˵��,� �X��Nutθ���lw�0:O~n�������n1+?�i9�h��Q=V������B�me�BA��bdxx��p�	d�`ߋข��m�J�~��\�w�q��.jJ��� ��ms��������������<�G�;���QU9t��ݢ����Q�{��$��e���n��w�	�E�\�t�&�p�\��D�Մ����l����8R��j��zC2N�Ć;l�������IH
xV��>S�;���X��d`0j��\v���� ʗ��n�O�n7�LAU��x:k�����i��Re�ot�.�L��B��@�:Q��b��q���CKn\�=�Ac�D	+�v9���4��l
x�U�Vט�$a����t���5	
x_���ǉ6�Mf�Ӵ���3������ߺuKp�"R;g��1
;�i�8�Դ�����a:��`�Y��og_����65��eo�y&���BJJ��$�ኇc�jF|k�a�ϐ��8���3��rW;ށ"H�Ծ#�A����u�E�;w�|��3ߧN���o��	�4lڵ\�	�OL<��U�E)I:ن?������,8HKK{[���!GѡX���љ1j�\�����@���m�q�n��л�Y?Ֆ��:��o��)>YPHH���fB�CK�8���Б����ˆ%=��I�^�X�h>�t������m�lm-�7�J���yo���u&�o����M�y�������<���<.p�5�ß̢��Wf�y��`�ǐo�m`9�p.������D�@��-R���ֈ{H\��إ�Lw4�\�-��d�[ԩ���.5��J�aH!�`_�ĩ�|m�S�r�I�,!!!a���j�O�!�7��kZ�Զ���'Vu��f+�c�
��I�� �ށd�U���z���g#��=�!
Yz؜Scgc�7,l��2[�+~j�!�7JP�m�uc@�!p�z�!���\h���%{f�QT��a۠g�efզ�ׯ_z)�{6�x�,0���BB:w�+��G�����o��h�sj%:R=��M:-�VQ���v�T�-�u���t��A�����ϣ�[z�W�^L�;��w; $n�f\RT��#��',��|q*P�`dQ�r�~WTh�:Ȧ� ��`����a����ʘ�����57b�¬Q�R�t"
5��� B�y�۵�* pr�)�AH�r��s�#:�����t�VdED<E����8����u�vC�̍ݽ$і%]��q$frz�C[Ձ8��E8����ѽ��
Ix��:��O�SĽ-�"�:=�@+����>z$K����z�sT�P�=����?����7���)�W���q��l�3����iii�jeG�<yr�c�=�������د��*S�y�?]Ȼ�e�1ӛ+�Un�؍e���~�~��u�>#1 �ʆ�t��i���qٟ��������}ͳ'$$d,�q7��hD�!|9������&�+���E[�v+Mj_!"�G��G�n���p	k�jk[�0[��#_�J/h*�{t�g�6�M^^��b_n�;J�[$��*= �u,�쯞=^�*j�XH��l��{�E��lV��>K��JX�6�Iq��R���{!@j���dh�y�`�yk�l��-��9G'�q�M��J &y��*q����E9�xI]]ݗS�	���i��850���G}�Ap������Y��k�/�WCX|�=�_�}�"
���,�����y�}~]��,53ߩt}{�<3�Y Ƴ��#t��A���,)t���AG]mlX���û0��t݁y�h�^>��Jy빔��`ɯ3���馦�PYIt� J̏?*�N�s˂%�f;��A�k���Quuu�dBCty����'wsU@� 2d�=x��_g����!W
!�����"���E������X������o/RǨ>ܕ����n��AA4篋�E�@H��χ�E�-�^ۯ���m�o��[.�D������b�f}0Ͽy�w����1�	��S�o��λzno�R.@Sz��K'$$|�
��.[<+���i6^�戳�	K��� xI]`-tuE�#/���J�3r���n�X��"��kSr{��I�ݲh���S/A�.�0�8t�Z�h҂�\�ל�@ ���+�;����>�����
�}�Ǐ�+ʋ|�Wj���B'm1��f�Ny��ո�̕YT�k1Ĳ�AZ�Ha�XrN�/�ς���~��_e�Ҁ8���j$58N���53��Nh��S-�󂘴���sA�z<j�/K�¸i ��ꏇ@���D��� �4�i�����1�����

����� b	�7������5TM�.��e_�+әλ���An�577w����=|���OBs�� �Y���\ϐ5�c�&��#.ct�7�����a��=P�g�cw�:Å�������lb�����!RQ�����;��Z�O1f��F@�e���ht��ۣ��;����~�������"�Y�s����Em9A�S1r��j!2%<�H#�&@L�I<<�6����U[���5����s��F��C����;���(��9����c�>ѡ�%@f�;��k0��!!YLe�'ͫ;�ԩ�wsS$:�܏n������m,dgg��*�Hp��(�I�'y�k+�-�u�fO)���\[��w�6x���N)w�=�.1���ʿ�O��>����o',i�[
(�DWo�r���]�hw���������]$"��}���˭���k=j�t'�v߻rE��'�k�Ĝ9gǖ]щn�{Z��{�x��BŴ�M�^{���׃hG�$�_��|���f��>�����ü�h�� ��X ��=��y�����O�8�@�&�bu����с�>S#�����n�S���A,ӫ��h�E�\�&��S �k���-�a�
ہ�{�W���a�|�S�F G!n�t��.?Rt�����|�F���O�hg|��������eof�wJ��s��[�A��6-���R�Ac��T�k�~j�S00H�� ����"�,��{ ��ƅ������ix��? ���3Eװ��.s<�Ob����Ak�j7�Q4q���8]��|��5�r[/� f��P���� �U�V}B� ^�KRV�����Bz�P	�MF�3�����������>i99!mqQQ/��7��r��[���o[�4Q���d`�-�w_Yo���JУ֨	���`��M�<V>�L��
���'��r!�:~�������ԡ��&:�� 5���˪���-��������������L�x�y������pϝ������G�zċ-��w����^]]]���������Τ�����L�����/0��4��E��\�KU�"?��浪0Z�i��p��
)E[S߿�b��L��=F?n��{�G�K��Ʒ�Ӎ�z#�Ή��.�	1��Q��G���?��R7�|)�A&����h@#�9��+��ཛྷ�Lѝ�_b�*Ĩ�&^<�],���\�vG�R��"��9glL��vQ���&?I���$��AL�7���C�+���R΀�����Ni{�B�z��5�.۬���v������#�i80��m�UQt���Ǐ��N��"t���)H���&ZH�%S>�+�G�w��w�T�����\��ߴ+�y<�$D *�s�2l���^9�����"3���>0+�`C"!$��j�����K>t9��s��Bب+S��qH�B�^���c3��ݑ���2S"�#�߳������@�4�c�����?��R��O.�NK�"��jJ�u66���atAAA��*f��� ~c����yÍ�ˇ:U/�?64LQ|�&E`�0:ח�V;�I��deeU�^����)�6��:u�����^�N�PάA�����5��+� 1+]N�f29���ﮃv�����f�E�*R�������uI�@�޳�4��{IЉ��|�)����C�
���6.]��)i#
�K����R\b��J�S#R��O<-H);Kߞ��lqQ�)�4�S6.�etر��"6��_�t^�Y�m��C��ڬ�H ��9�4�R?���
�,�#�?�w�'ɺ��6�oN)���_�>�؁Z���_v�o�Y����c2]Ml�;�G�C-�Σv�m#��gd�W����O�x�����`�7)*7K�x�]|��L�l	�������,�b�LxCP)��>ˑj3����썩���NQ��O����(�S7M��B��;��~W����бj�!�R8ۥY��$�x���N9 G����ɣo���R��,N�5qX�P�����V鵙N>�B����4`˼�O!���SG5�-u�e	�[q��cЯ]���o�y������(�(��}��2������\�rV��jA�������C�����;�;�,Cn����8���ħ7�,��ׯ��?�#ɸ,*])��6M+�=��Wz��:����V2���xgP[Mm(��ε��}�����1,�g7	}!����? C����#��ͱ�$9�����U��C��E��Ԓ�����&����������Ι�����⵻�.��9�0G���&N����[��堗գ����M�������SE]�H�e*k�~ ]qz��r�]�V��gE��NO�����܇---|	))ʨ��63D��{n#$T�866f��u�r�:^���ޣ$����8YV�YVl�|
�,���ۯH$|�:�(�Zw������8<>�Tw��5���C�H��p��q�NGW������h�[�9�^h�ziwޑ/j�r�ұZ��7����=k��j �ޣ��) �kڿ��F�d�~~��J*4�М������*v��=�^|�2ǰ��I��L$p���!�g�О6@֏T�n5�$ǼH٪�ɸ2�(��wdԯ�{����8K,�NuvʎG�;W��'D+�Ͱ��l]�Ұ?�Af#NX8�O��5N�ڕ�l��8�#�������7O�S覀^3��{���O�6m�Y��N-��`F�������G�k�Zr��s`�A��rZ��O�O�tɷ�/F��W.��[[6AlFa�3���q�0|9u+���-Z(����r��6q���Va!��޳�O��m�|a7�4qħ�f����.>�TM�7��mȸW3��(�O���QI.&>^/~5��[��I���!{����I�E����5���QɃ�qog(`��U,	�W��jѻ���+��g�-f�ϓ7�>������n�h'���oO�����䪕��F�xl�*=I����й����0��>�l��6�j7�RAW�"V��
��Bvz��J3jAgBXL7qx��MJɻ%"u8�Ef������b��UI�(�Ɠ/bZ�9@T�.�<�}�����;��q:�,����/�|�!�h�����T��=R���Vٔ��.�m
�������9���O�tA|�����Y��l�2k7����˹�;���j�W��Y���Td�\o�^���t���Sj�[�X����CF��3�Fd�f�/Kș��S��&>g�tw��؝�,4�uꗑ���d:��a�D���| L����;4YE&��l���P������č�����SV�����~]2V�C�r����UaḶ��5ytS�v�3s%L�o.�u�s�HI��}��jЍ_Ihm}nj���Q�X(��Yrن��K }}}���eV��ܯ�u���w�{y�����^�ǻu��������;�m6~ݺ	)�|U�{p۽�Ұ������"�;��^9�}�ȹ�/�E5�(���0�7��M�rN�1<�2��7�t��C��]2\��D�� �4��_�-{w"���ދ�?k�!�����A--��Dk��w��0��9�抇q˩��e7��6��u�n�h�hˁ��0rX&mko[>ߒ0�/iz���/�Pqص��	�n����ffC�f�'' &R,��
����z̴e�q	\;5�F��\���'��;�������R���\���3�Qߔ0f����)�/Gv�5�b�~���1r�+��/�D��X��m�gӨ�!V4.����.�ё���Ϸ��o�t��%N4c�[5�>u鎪��̕�_n�����C3�<k�e[��� '��m���{fJ����r��ŶbjGR�d��۷�ֺ0����9�ž|uqq1�_Ev(k������d���z��gބ��T�����!�����t�|(���;���b�ݣ�����*P+��%#/��Ub�3-z��v
1�Ą��d����8�~�� I��~����fm�������[|ލ= ����w��J����M^���w��Lr_��H�TT�oN��/����5��S��ᆯ��bk����1k�_V�����֨��C����������pǢ���^*Jʕ�����\�TЃ1�5C�ܙF�@��߶m�����54b�[Z�Z�X��_����1,��T�|ߒ�w8�>�����P�5aA��[#�A��OnUV>Aߝ7Қ$��q�L��?
ZfY�S�i���w�1'���N _��<6;� �&��#�Fd J�Wc?����gϚ��K�|�����!@�s�t�v2���.�$�C$�!XJTB�{Q�F�AH\\FW7�@���t��YO��u�9ԑ�g>�bZ�&���H�|Vu{.f��Aw�f!�E�(��L�����{G��e��S^M�W�Z�x�x���6k�7ANDDD9)&��BI�A�m!i��"������YL���ѣ	t�L��7��[׮�4�B[��8?�x�[��c�`����lr�(�����ժ�*�(oR6C5]]��"� ~R!l�4�����2��4��@/��U��M��cp�q��=�K���	{��=�x��А��=3E���m�/�0&Bs��Y-�c���T�z�mv=t�b�\�&��K�d+>w����01V��Fw'#y�DP4��#�������Ы23��L
�q�B�2�F�zNv=���TW��Kȭ�M3p������{�9�/�Ys�'�+*�Eg�����^ZZ"�t)��ڜ0@���o�V��#��n��G��c7�hk��%��N�u���X� �e�>@����0LE��Z����w]ؘ9������|Q�L�18�}U�c�|�ɴ
r�6#lz���LLL�v�zBXƟWكԻm�9bw`_JD�3�I�f��z�-2˴���śuF�,Z���.1�t��7�C�ߔ�y��7"��_t~��֗��wúg�@W�ʤ��R �+�W<6::�>�aT�3�`6Pd��1�:۳����߼��)��>o�ru�O�Ag�&f
"�a��S11�0��8I;�MLL4¿�}s�΢�<Ŕme��,��\c�9��d��Vܼ�E�z�A��iih��Hz0�V�U �ꬁ8�A7+7y0i?d�ܙ���]7kmm��m�����]�Ŷ=�+41�7�ͥ�	*A�)�qv���}ċ�}`��ϟ;s����{d� ;�~�Cv�Q����t�-۰/mi�4�V.+H�U�jȹ������VJN.hƘ}���|���>'�#_{}�o��\�r�EN��^%k�g躼��d��y˙N� e�������x�Be@�Ǐ�H�J�&o����[zO�m"x�le��lD���C|?��>K6�ثvsq!����e�e���f:?�nB�		K��$�`t�kF*4�M��"�h+�#�?��4����F@�0�d|�fuc�G��.�U�(9���t#V��'�>]�ll2 �<�1G�Q�b���_�t�c��1�\v�o/R�����R`*��nT�P��t-'0�kO���� 9��|��ed��o��F�;8VVUјC�(f�����KjT �:����b�	��|cA�EB����vڗ/�YXYu+?\��BS���O�����o�J�Z�l,��L���n�v� �<߿�f�zu����X�&�#$:�0��&�C�y`�Cxh�]{�.�"�썌��Nڌ�Db�k��O�?��!����A�q=��{��3���5��!��q2���4������RQIE=d��uG����1] %M�����qX��=V�������v���5�մ92]����Acv��1Ϡ�n��ppp��*�+�����a�v��,T����Ң`
�=��M&��<~߇�ݙ:ѣ�/!�{�3��$%?��wF ���R��s�+y�L��8�Ç�-&;B=�T���|�>�5�"?�GE;S�ײ�&� �>w�\���Ͼ���ݱ��5c �8{_c�����Wۦ#7-M
m�ە,�be����Ĩ���m���ʇ*��$+:�c��S�j�M�zF�VK��Yn�����pf!Ǯ�	��}�j�l>�Х|�QR�'V�0�������{�2!�}҅������w�8/��$^��	 ��b��3���tz�cJ��������]޽�Y�h�e	�h<}�N����H��3�� ����i98���^�o.�h��Iz._�EC؋S�N(�i�~����w�����J� ��ö�?�������BN�S�)��y�A��{�| Jm�>����B���0�q��c�?F7=h�k���#�T���
V������X��F�ߞlj��;@�r��=������Q_Skk�+����~��emN��|��i�� ��"/�&-mH.�\G<��ȟ?��@[qqq9�"�)��Mg���D�nMRդK�k������H��|��vD{vz�﹖�mY�7�z F�X[��䙚�β��?P/͉��g���!!��=/�R��W%ϕS�g5�����\��W��5=���6.��yz�]�O�����p��33�,
v�t�r2���O7�����)`h��wb�SOOb�|�̳=��~�.�vc������ɛ�,�k��Z�b6>��E�Ƀ�A:��^�b�5�e������w���zv ��7��oM��z#`B�GrP���b����q������.r��Bc��������-8C��B�Py�.?|P޻w�<�Vނ���;,n��4uk�'0	0�7oݪ�n�'!#��b.%���y	w�nA���+�{z2�U�����������_��g]�p!����~��p�4!!�+n�=M�ByԘ���߿��!�S��f�"�6C�.���aQ��?��4�.f���Jy���ge��Y>��z��&�A���8�{��'ǨÛ�K�3�
#�ۇ"�C�V�i�Ȇ3|�����]�~�C��#��Ds���jH�v >�@Ȣ�NbR����ײ����#����y�S;B �o�$i��<|�0�a�K���
#o��f�9�q]�.��֯���r��(���l��y�Z�s9���鎤����nolK8v~ ��u���lq#G<��f�t��=|HJJJ�z�A_MC��� v4��#ᵳ�65]"_b���1羱�a_?Uօ�AjT_��j�Y�'�YS .��Y3���c��%ӫ�]��~h]\CC�����"e}Nl�4<��|���hrz�<i�gV+;�r�0�7�o!b��k���rN�S���˫�:@1J�>��� ��[���Z�����!�9�^ �[uz����ڜ3T�q]+����Jt�e�S,6u/Ş�L�gߔ�����{e�������	�8q��wϱ7B�#�O��J��TTԫ��\9� r���c܂��
�:-S`������:�ۋЊ�>kh�9O���G?�@��y�O���Hv&���E6/�n*O��e���T�����$$	:-qHM�a�KJ��W��&x
�����9a����-&��S����� ��Q ��j������E�����?J�hl�����],�?Ɏu�����`�BS��t!(���4~GW#�kR>��.�.��0@p+>���B��&�$������o/Q�}��\bųdd}�1Ԥ�����2�y2E;�'��u�̫��������ׇ~���߂]n����"nk±��o�����i�~������˫�ys��\�]u�����'�)[[[�a��R�f�^?�]񽲲��?���2� 8�C���_C>q%(L���t�{���{�@rq]�`0�
- j�>�`��;�L�3��G�\�o�#�ᅡr�=�^V�Kѵj��e4�kЕ���Y:��]�;1!A�h�	�4x�6`~��$�t[k��[�n=���a�5����">��@ [lL�e��r�X�-֍��FθFצ{�S!It��3"22�l�
�<���x���������8o����i/@V��5S��6BS���C��8/��������*CT���z�=/��Bۜ��tY�Iכ?��񩈆�N��� ���������ӊ�`��J�(�(�MP���q>|�t]}�ܤXBW7���o?~l��ի)���!/�Ӱ��r2�������Ѓp���v�!�0}�P�En=J��G4�Y���ν���gZ��+(�����Y���B�9�x��H��j�H~No�xI$��}ȓ��	�>��\�����"R22�SI�{>�L���� e��̷�VWW�K=}���-���D$D?�r!�W���Sc��)\R����	����aL^�N�{'�o꽍�v|��T�-&��m�ޑ��!���o-�F�E���0���"��"{[�$4��;��&��j�3����Eb����J+ڗr�@�f�z� ���qT��_�~m����M�_q�Vx�\AFF���E�ǥK��0���������0�2Yk?��q�'h��#=@�Ƥ��6�..�� �����"E�����8&#5r�Q��u`��M����L�q��-�������-S;W��P�l+���f�c�7�����5#�|��q0��@p�{k96���/����@�X/�x��<��1��/_���vA^bտ���#㳿H��=�ʞ*�&椭��+%Ĝ�����k	��/M #�ܞ�|SV^�3000�@}{�3�+�4N����77���}��ԋ�~k�Zգ���˗/3�8������Qw|N?H�����BCA0�9t5zr�ӫ�B��C�M8C��\�v�l���)�G�@����i���j���j~��~���-)��}�vE�[�>��.�Jw~8��i�wH�@o��-����x�Wܰ㔁�!�sș�s�t;�+In3qU,�$�K�8Pl�+ݎ��I�d~+� �g�8�; @�&P��E>� �����X��Zn��3����B�
J���������QQ @�II}��#��{"(�U���R��]�c78.{K>�8.���177wk���認� ����_�%��?l�i��>���\��11?��1�F���"ǵ�-�Y�J-��	�8edA�rJ�NQf?$����7���t9�81=������y�vj�W�<#�ٵ*	10ys��֮�&���;{y��aAhv�潧f�}�h'�\�`.����(�r݌�ׯ��0*�R�>��'�ĵ���n�La���d��Cs��7sB��;��e�ߥ*���y�����U�X�);�~�|���Ғ��Y���c=�:�
��>�[t�qq��`��+z��]tF+?
	g\%�l���{r�=�������u��Ew��}�0w�����]�U�)E�T��6���M�}=Z���#z{C�M�bM�����z#do_�3Z�'��Mƣe���h��]NK**~�d��9��d���Nm|>�O����Z�}�ϋsG*�[$����/�Yf�Tm�!�� $&�6��S9�縿��0�	�+E6���\���4u�,���l-�PN��#����zH ��E^f=�d�MÙ�쪜'�6�:G���ʏV�b��P�g�NA vrȕ"[��������3{���-@��ڄ�_/���Q�n��&>9�,hwq�C�X��G^^&��ꊪ��̌~�\���-F��-�E>*ݓ���ʨ�g�
`cW�?#�zYS���@o�`���{y_���?�(��{�Z[Ay<9����5o؝V��USSSUg5*�c0�k�x`�۾������k�|9v>Þ�n��N��N�ᱼ�<:���+`�� ��p��^��y�N:٬>�+�g��&=�q�~�w�s%$U���\��=F�}���܋��!Ă�V���$�W����8���rj��^��(@����K#���g�\�OmPX�1�\���S�K��F3 �	 ]iJ�
,�ҷǲ���X��a�H�i w�Gj��X��?�q�Nbjjس�ϟ��<�a2��>M��\PP�.�-M] )��x�$�ޯt:� o,?�V������n�^ݓ�1�c֨&<ik�-���6k�->��,:}/��g�br�N��f��SBv��ڭhE�/�R��;��kU�Uu��[9x�<�:�{?��i��t��%��94Ԁ�?��`��WEE�7�w��l�Ll� ���n>�Y�*z]+a��3�ߚ����c!�e��?�7�.Ow�jxP.y_�B�+%�%�ה1Tz��6�g>�o7���%�~ۂ�3������Q{w�|����=��7�6ߣo�XT?��I3�N��_>1h�d��6�~{-N�Je���fՑ��F��gIIkԹ��3���Ï�oMU�2q�E�� A����C�T9��xS�$+�$&&V�vz��%���I����B�ZgT��Xs�	���%�5ҡ:1|�Z�kyd|�M�Z'a|�i�|�d��ǎ�,�����_o���6̲|��d���W�Fo��
'ɤ�������c
&0((AIuM�'�	m�����zteh%!�ya�Pz� �T1�U�P��� 
h6g�p[�0�nפ������ʤ<71I�dw�����3-X��O��.��^�L��*�%O �7��S��Z�TT�8�8]
�&a��d���1l9(��8��c9�@�袓�v�R~��	x=��l�z ��"�c��ɜ���M�k�!W]_�τ��-&��t:a�b����W��l�9� R������i��D�e��.�]ڒ�5���JBLb�W�t8�it�����i/�O�<	O`����SZ�oOS�jɎ�vzõ�.�D1�]���)H�Ʃ�$�W|����@0e�r<6+�?LF��� ��ԝ�t%Ԙl6�c�Gh�akڑOyy��r��~5c�yߕ�OUIE����v�˙W��IC��6M5��j�W���0+<|�f��q�! :̋65�|�9Ş?�S2��C44�1zP*���}�'w�/مl���L4^E�kk_�x�@R�����c_�o4�|�^)�@BZ�
ô����*�ʀ�oIר��N/��+Y1��I���d+�?hq�nFdȚc��X��]_0�zXK*q��&���~���������� 8@`��6���G��1��\JJgw���#��zY�=Й��y�fa��pH��ˮk��~04���qT�t|�!=���>g���`���^֫iiT��u�6�1vu�Q�5����3�F��Q[%R��6~	������/O��] �^��x�+$$��МX�����G�s�"AR`2�O�av�$���]L�/ׅu�(qq\>���W�7�Z��Ł9��>4	ld���#n���ʅ�UUUy;K5`i48�-x�021I=}Z����]Ů�b��䋒��/t�;M^�Qkk�M..������3N�={qө��2J��2��߽��Z�DKv��/rb0�D�TX��/��ho�����]��oI`5������|�3�E��	i�݂��0�r�KKKϟ>�Xn�S	P� yl��Υ���]���:d�9����`�@(C��UZ��c8��u��в��ra��>j�F��U��V?�w���V˅������Қ���޽�]{�ϲ��B�@P�hjv�+`���abZ]/���)��k�Lj�z'!;[����
M6��㨟Z���eO���o0%]�h�a�� ������ˁ��߇Y���&k���01�d��Td���7<�����`jz�sP�u�vm(��|�|�G�M��ƨ9�<ev�I|���ɖ1��3���eee"''�ە.����v�^*)�H�>��y��u���ۊC��y6�{3{8��������æ׿K�z��$&��,ۿc��U߶,��7�@*��{YĄ�F,�bϟ���9��#oa&`H�
��%!��3&��"iL����q�����r-���X�P�B �e(����@�"ۮBW���Ft�m� ;�P����u����
����kq����:��B�:�=#���u9��L9C�%�¸h̽�,]�q�ӧ�n�>��8�Y ���ѯwS-�>�##��n���/��.ށ?�M���t��]@Ω��t��nwƀLF���'Y�C�Fv��c��B�qw5o�^0-x{t/�zo��������]2��0�x(AQg=z���D"'��U�ڈ7o���]�j4P�>���I�3�I��o�
8#Zq���QyO9�]���"ϝ;g���8A���r�N;�A�8l��(6ha����$���L6��(Յ��+��J�߱P`�����zcނ̧��S"�`S�i<�D�?�nF@D��Ny8���nMw�~[����T��:�"P�9:��ϟ���f��GN�݉�復����iK�a@����h(�[=_��  '�`)�32V�w�����)�.n��o��;"�a<���72c"��+���0l�?�M�)C�m�ey��M��W����s��l)R�h���컛?�o¨�r�'��˫L�luU�&�1++���AFL�LO7V���xC8�V a�?YF�h- ���J�x�B�\�jN�^G5�]է�7��1%]������h�ې������D�Ċx�?�}��1.:ҹ��mr���������~xX�Е���D�TeT�洜���se�"�����?��w�N-*RF�6����H�G��T>���0�� J��1�7aJ����j�1@����o��^��+A>
����L2��f]��u��3�"�1T�x@[���F�c�9AdL�5�7��>a���+*~{{
�_WW���f9�����k�lv���,�&J�X�@Z�k]Zq�%w���IT���CK��:# ���IO��U��xbR�����3��˧JpG���[l�8Xc�oG�&9�b��5�1}ή�����>�<�Yz2�I�U��W��'�6t���0���@ ;�2�)7d��m���qbع�Z�nB��j�-�>2����kws	�孪�%����5��������|2'RRR`��vFo�I����zp��o.��~��ll�]�X|ލ{��Qwƛ'��#�)�%@�f�GF��_�4%�%��T	`��k *���k�&��v��?�TAGq?�)\r]�݇�ld�;Ñ�^qT%��\]���r���uoN��� ��{5�����aff�2�	�,��9����=:�c��`F���7�Ο��ucêeQ�BM�se唲���
�5��q1Xz5���eq�(������X�V����;�T6�����[PI)i�ͱ �CS��o���cΐqVzw�~��) �;}��q)V��◢��1���h�X�<AEӡw��Qu\����E�h�S��>�v���{E-*ƨ��L�	�;��N^Ĝ}�`<���>0IУsh-F}�R���ETt���)N��[44�A��[9ur�8'��*	11�TVl`a9�Bњp^�>�:�#����g�0����g0vI���24�g�2D�0ᨵu���y*~�ƥ10~ �a�4��G;��8J\x�O+R�� ��@tc朧�O]��@:ԉ�M�s)Z"c��?�&�! �pqq}c���Z4�abQ5�֭j�'|&SX)�`�1@�>+�ژ�)�=�o������-�������g�+� ����jo+�c���N����$x^ggg`1�k�'j5�)c�[U�ٖ���V� �|}���������|(hT�rŧ���]X0F	o�`"��1ȋ�"S
^^^hi&-WW��X��8��St��8<��NwZ�!B��i���s��(��s[�#����,���򟺖`=�'�3���R>k�s�� .���HFu�56`2�@ZN 0��Ł.���U���L�h�� 1�� 6�����sNE6Q�ϞEA跄��J��{�⅘�#�nH@@p��#_M��i.��2����T62m�p�pG�W,�"��o�k|���!$*������+.���\\t	�κ�~�%	���M<��f26����rˬ/�UKk�$Rp�>�D�k�x
ђ�����ߤF�d8�����p�-������MV�5�bN�-�q�(�yM9������q%����K���-��J�6��*���ƶ������!��$$	nn�Q�t�g��v��l�с�ί����W �ӧO�/J������y�v��lbR�A�4:�K�j�x�A� q�
���^b��;@r��8����!R��0CΓ;N�C������P�����|!�4x������ory��9t6�޽{7��c�������0ڝ���	C�%�����?q�C����m��"�{ ����;
٥�}s-J�F��(AÁ�I[���Z�A)�  2�	{RdLՐq�y�ÕS�On����א��g�^�]��o�?���D�xX��㶂�@�VC���g��-���5t���g�ug�s��tj�|��1�*��)�
t̓�o6'İN ��3֌�r��B���_�0�wqXxKq��ݴ.3��O�]9��|dq����?���w4���Vl��؄̂���^�N��2oֲ�3�R0݅ͮ__��g�.���3Ja))�F������m]�S�q�-�Q?��G���elV&���A����l�:%C��TR� �aԨ&D�n~
Êd@Q���i7^�]�q�K�,��4��˟�� ��w�#;�~����T@>HP&��ER�a�b-*�[JZ����w�cu�顰?]Zro�A+�D#���l�@�V��&�Q�_T5����l�D����?��dE4LZ�~-U
�EL�%u�8ήv����lيs,�^�X��ฝ���1��(ir{j���?]O �o�n��*���`ǀ�p~�E�%xY�:�I������!��WHE�d�H�����+�����Ә0�=����[7�T�N�Κ-j�^M���F��b�z���V��xD��*X� `b3���у�s<������!���0r�&��2��7P^ݜ��ՠ�Ê����R�ʜ�.��N�}�� ��6E���@g�� ��5HK؋��0�X����9�N�Y��RG����i;�z�����X�'	Ө��9����Bt��3� �!!X�6�{4��9�}��t`H���ف�be�U��#oy�:m4<��z4��g��,��į7���vr�/8�`�Ss�מz}:%���B��)Z`��k����ڵGfj�����Eh�����X_�4�A��+�jos|����da>��B�b͸�����4+�Aa��M�nf����jw��kt2<j7��7V�^RC[XXc�gj�®6]�Zf�l���	�f�l�t���ק���K^���C�����՞Z@j���N� �����r���Lj����7�x~��F0�_4����'�Р�<}���G���FI���o�`k}�h[S�c4�(F0�͈��4)@�A�o����Cmq�A�4�S�a��|�.ƶ�v��ƃ�`<�����Rr�����if �[���ؘxЍz3�i���y�I�B��,S�u��wh?��f=�:��*v444�Gm����M���;j��X^M=wvqٺ���ݽy��/��ж�3'2�p }֫����)���1���܀�)���8�~��
����(�>������0�п<���+�Y��M�.T���ؗco!"≚��&��.�-��H�fGߞ��!J�u�i3 ��.�OeUe_c{&��F�wv�)��� �x�ʬ��x�zD��P��_�Iw����`o,��z��uT�E����jPoss3�I�[\3�[׮��c�%/f`kg�!d�[}��5Z���=��
ρZ���ͨ#�5���K��E�?�8�c�U�z)��/��Y�� .��kj�,��tt�U�{0��Ǎ���SiG���R�BN��***� ��w�n,cm���g�1s8m�o=>������dd��hCOp�\�Q|�O���"ݎ����f��Y̕����ޕ�5u-�[��U�Z�,`@AD��,�(hĲ��QE	�@���J�u�TR�%��U��f �[��%�@ț�������{���'ܐ9��9���f�̙�G�j�`���>u���#���˗Q��כt����|
�0B����d��� �{3:z�x����p�`w���B�aFF�m/u��Q�L2�n٩ �ş/T1|��� �!�R?r�05�Bn��F#���0Y�d��g��9��,Y�X���.�T4ڲ��rL۶��eVnIE�������1l�ʓ;}}C����a�v�.hَ�R��p�o��A��;r-�Kzp"^�Ԛ�1��UGk�:��Uj ���U,(��
�P9˩���ASOo
a�/QGk�v����h&���4j���r�.n\=9�ȫ1�u�q�+ 	��D����>0׀.A���W� �Tu?)	e���,/�F��09��
l1��>�����*�m��P��T�EaR��b���'����;����؍�(g.��'ǗO�k��	�5""�.*��	�S2Aɣ�Z � �I�S�Ĭ,ë�7P�.�z�y�X�J�;p�DRǚ�����Tj����%��m���d9�0b`���K������H	�(m{��+���a
"�6�7@�V0p�]w�J:x$�s;�����^;1L��b@���z_0&���=S\�T���`�+��~}i]ޞ`og�����w�yS��?�(��?�������O,��ٓ��\q�ZzNsN$�ơ�n��>��6��lcS@؅�ya��'WU7��;�"��XH��&!!��%h�$(tr!-��ח���b0�R���6��V*h<d�����M���q�el��R8k�����S��ibt,�I����vD[`n˹�7� ��A,�8���x{��`�?��o|d�S,�IիJ��s4i�K�MiPY���u��[���5�̞w������������e=�^A����{���,��\eu�xP�nU\�EFFF8�� �C����i�9�՗_&t�cu�I���B�Oo�XS�_�9��'���!��B��ҭ�we�"Y��U	
<*�R�R����ƺB���OiS))hЩ�F-�}���tk�g�d���~����ǌiow�A"��~LEE�����&��dQϪ��<@8�ɻ{`D����Z�5���Yb.��(�u�nғ	y�P4�Qkk���\Lv^FY�h���g�A��}����n(�i25	�c�Fj ��"�8��"o�@�k�6�ڼ���O��o���N(^��12Ŧ�}1 ��-#k*1
���3�=8Ҟ6�.B1/����L*\��&����?^�R�lHƚ���^G��#%֥�z���>;�V�o�y�ui��$����Q呾2�MA#T�ڧ��Т�k�?���_?~���g�Ș�\�����m�2�;�	��P���K��IjlJ1A�som^�9�5ľ���k����@��Mks�����y Hd�~��4���QzM��K���c�>jn�: 9�<���we%tq����Ͼ��+ 6w�G{x�oJaJU����Nk��D(��Y;��jc���[���I���\jA�X�=j���w�;�|�����t ��;	�4��1�o�U������q)��[\aEY�G7S�-^��<�0l{ɳŅX�V13�C^�<&��w��Uk`�0���~E;�"��F��><�������<~,�s �3Op=����b_V�.5v�f�vRo^[<�itHd�/���*�_�e�h�YE�6Q\�|�^I�R�ֽ��3ؠ�>]�
`.�W}1N�٨��;�4tg�"�1�;�z���e��{����P$V_?GBA;��Դ����=�z��k���*�~�m��e:5�t���O>L��upw*Ʈ�WB�����$4	pm\�լ�^#ŗ��f�)��f���S�(�M.���Ӡ�߉�[Z�r�xG�w���;���3O�i�Y�����K��]��u�w�Y�7�c�#��r�X]v�!����C�w�h� WdS�4���A�-��`T�';:J>�W������m�A%�^|@ި�n�g_����fNY��^�-�xy
ѧ�$��Rmm=�z���� ��Ͻ����T��p�d�&��B�S�W�D�B����0�Ca����0x�SG����О�E[�6P���ѩC������ S�=��`��-X��`_[(���m���
˹\{N�7����4.�[g����/�1D�z��ؙ���9�u,n���m0��������8o ��K:k�7?}�i���2��?Er�V����wT`���B�����62pR�\$;��į�����i4ư��"��A��|��ja3�ܸ�y��,��8�Lv�͍d^��RQ��T&��zL+t�Q5|����o�ս�8!��m���̉���۫������qd3^�=5��;M���o����8�3���ߙ#�x����J�ĩ
��#����]�^򧕵&��n�ΙN�a�z��Y.�rb`آm� aC=>2_�rc�G:��w�"URω��*�I�@J6|@1L��b#��Þ�O��Š��Rf<#���`6��"�ӕԷd�+�$���èQ0V����|ڤB\��V��
f?+p��v����/�8=w�n��"��]��B��!®�d#�`:�+-e��FZ&��`v��6W||����)��@��EVJ5�R����x�ӂ\{Ir�i��ɓ/�G��0�4��7���l���ޗ\���8NNN�n�v��Zo���N|�3g<�N3XWu����γB�cVff�����K�>��ǚ�%����>-�osQN('��	�rB9��PN('��	�rB9�H8X�y�|��6���go�)�����ˣ����w�p�2�љ�����>�7�M���B������?0���C3Ev�u��f���r�@o���A=�$hd���E����������f���]�t�����ak������PK   �v�X� ���� 
� /   images/38cb4f51-bc72-4d24-b782-e5d855ce8001.png�|gX[n�c��"D���  M����t)���!�H�.���*��@@�tB(�	�����{�ϛ�<<g�^�]k�k���*�2�etMQAV�R	���"�˅�_������>��B Ǘ�*@@ �o�/Q���&�#���sGM�׎�/�MA���|�6�&/ߚ��ڛŭIЁ@�@���\�W&\]L��{Tw��_����(���i�m���?t]l���c���c}y0�"r��n>�~�2�4�܇���y���:]=�*���u:�����,V�;S8ܘ��`��������Q�x�_���YL�F���N�I���[̪��9���?-�%O�I��;�rv(Y�J�ӣ��7ǉN9.]^;sn���g��/~���7��w�矤��2�Oߒ�~f�s���&�`O�V��2������[�
�β�G�~�z,�x�T\�Bgv=�@�(��5������ЅM�9���<�T)V��m���q�X�
k����8k~Y�֖���Q=�AٗmYo� "�~A!�����K���WS���>�7��eO�r�D�ơW!ԁ����F�{�v�ٺI��G��h0ՙ]8jY����o�/8�\����q*���⩛6�萕t��嶋�Q��E����Ma��?|)�?�晬BuGQ¡S�wf0�'����򇞨�����?�����}oy�{x*��h����,���B�4�*���caH���%u<�@�a��%���{��PZ|g�$Ӑv��+�>F
Z|�[\�U��5���:��Gac���|�{I�5�݁(������Y"��S�ʨ)^Q/��β��抖��h��/�Jq�U�_��:\�K��I��\�pk�*	(���t��Rj_k��i�z8-o6"���<7��f$Rv?��&hD�K�ean��AO������5[�U�tB��&�lb5�53$f��K_�S�j�nl�C[A ���>��fQ��b9���	Ysl��^�䟧E	���"]`i�ePybГ�O��ݛqo���XZ�GXP��؂�J_�]�Mq&(O���������O��oW��4����L���T$mW̄��-�-��w�
S���<��f��p��)k���N�j)����s��y&D Z��!��5�G�D#=�g��B�*�kb�^m{b�R����P�xs�s=����� ���R^�j��)���h+�ݰ����oF��3q���#��W�Ev?��b#�Ќ�C^�,�U�4����2��A<�z!�P"Aѓ]���~#)Pz�:q���Z�z����A��Un���@W4������AK�WI��=�5���r@�+J�:e/_��&iК@om��*�2h��w�0*��;7(�#"p��{�갥LƇ����	ý�b����W���ވ��DA�?)^�k�d�\X0��;0�FM2�%/�u���go���ܖ�Yo�� BH B$�2E��o;���v�_9z�To��yK�b�mFrv����f��J ̴(CN�w-�)�zܞ�1�i�Z�3�i����Jl�Y�@,�Q�=�kI9�N:[�9Y�CznE=��ܓk�k]��l�q]G<�����T�D�P��@�[�I�қ̺��e|�������k����dr��r@�B��S�VIr%Պ:���B`�(�i���W�t@x�Dp�o�) ��jN���j���#��A�qN�U�8�cE�n68�S���3b�A�
;yTr�}�Ȏp�W�H,�j�b�#g3��)��`F/��qYh��i�/sD�/��kF)�h�4gy]h8�����q�Y��Mh&�$/)�j�7K�zpb�;˥�6��Q;���S�1�G<�?���ϣ I�I�4��t7����bn��:�q����6nDrvn�8�LVW=�0i�i�~��|�n'W�x<*�L�-2	6�eDZ�k���
c�@2�sŧ���#	.�X��c�X�;J����t�df�� �OS�U+��'�f��N�atn�ɒ�o"���
��Ū�A���"q�O�7z���5�:V}�>̐0�RB�@�
g����ӊ`2�9����L�fk@�R�wђ��B�z�_�04n";،K�N~�g��M-����?�?��8�Zo��U�~o��*yȩ�ʪ�#!���$���|I0f�g��
��[��W��s��t��a�rє��p��ӂ���a���z��ꅖ=��'`%�������^��2�	Z�)XKS��DS��U���LF��A��S�å�X�W�3����H���_�\�+x6�xN�3n&؃Z����Nշ08O|g�����L֪J����/~[0Th�r��T[���1�1�)?򥨧�D�RA��S�o
_�!Lv,���zk�21 ���~J_"�&�f�=S���Sw'�^�}�����lbm�ec	��=/�גU��T&�BK���+�t7���l��W��͡���D���,c
&]�=-����xUV̒� ��K�ˑ&0Wn��Ǖ��s ���*��� �f�I�$/�+p�{�T%�U��O]�&�d���i�\�yꉭ�9�-��"Zg	�*��dU-���Eh��oe'v�N
_��}d��g]0��c.~�R���H4_?�1sD����\EA'䢬�d�X=9�� g|�|��FDt�Q���6�B.ҥ:�w����ZZETyVͬ8��;:�s	0��hЋ����x��Q����8IR��<�Vv{t��Y?$�f���<�/
7���V���!D ��S�~�J�g[^����e/77 ����~�9��-�p��%!D	ܥ� �	FaYAwo��-��J1D6�	v�C�Ӓ�~�GP�(�m����W��m�rsr�S7#�MF��������yyy�ɋ�FjM��FK9˭�M��w'-SL�7B��_�/�.�<#��eRHG�8�(;� *h�B|��5g?���(�3�ȇ�'�;�8�>k0K
�L��1zI0���،��D�S�,O=F�;����T��-�9Z��n�]St�#�AB2��'��)ν����(S%��T���3M��k�U݋�5b�~VT�����4��e<4*%�\�㟣&,t��ds�ψ�]-�V0�r�����o�� �����SIb��Z�w��d������e�oie��bA���G̴�7>�=m_1�Y�yN�x����C٫��߿B����&�gP�<x4�
��OIIi��4�Xwk��u �<�W�_����C�-s��L�����xݣ�J>ս;��Vxhhcס7��v�N��������Q��L�ɿ"��٠$3'gGp��V��F�&Nl�-i��2,x�|w?i�6��v&D��S�O!hm���$�/|N=ӗف�ޤ$3�88 !\R'�j̀�K �L�">Q+�ZZN����1c3t��\}�������oIf�ۚeeeFIǎ�^;C�����!Bx���|Uz��P!�������%�*�ԙl����_���b�Ť?������1K1��f�f"����]�8�{�$��YW�K�aM$����C:�i�%!Ġ����n����ү]hi�Bլ�uBe)����w�rg��A����k��nP���ve�4w�.0WCU:cZ8����S�������inW�7���u����R�ʢRPd"'�;������ѯn��,�~�`Lf*����Ò7���
�n�l\`�GG���x��7=T��'�W�睘�S�q�B�ʥ�4�_^�5�E7����Y���0}�;r�C/v?�cY�5ag\��a��R(-T�4�������I���[k~�ͮ�<����a��I��Qx�����W!Vf>�{�mk����VlX���f��iz�K��x�x�ʣ;*��x2�t�����OK�� �뮥���N~d6	S<P>>;�3��!i��gj�5`�L�8��p���/:$!y�Fx��U�
�V�T�ZUB��F�w]�^�9��D� �OAqf�`����kג�����XN���f�Su��wW������N�� �#���z�wR�s�f���KC�ڿ��M3���z*���e�I"B�	"B�f�,�Sb�,�jsxHa���rJ����ؼ�^Kq�8\��>0�0��
�:̦x��`|q-! $·!��̨DO���_�R	�{	9��eſq6��b��܀��w�q����Ԗ��{��r(���a� C���M�Bk��y��Q��T�Z[�l�0�*�l;M��ٕii~^(�HY��<����n�0 n��U���@M�6!��$�_{�#2�8Z󃺑2K����6�R-�S #�h��s׹��cNqJa�q��]�q��@�2�� 3�.�\!ݽW
����T��^l�����8::�2�]\����u*��L&>�;u�{��zX`�����P������Ͷ��x�;ف|�V$�@}�ڲMq,3ǥ�ӓ���<�t�f�TދU��{�Lu�6Z��Fl�щ�&y[��V�_]=?�+�
��v����p�i��{�+�M-�h�.j�{���}�9���bO���z`D*��
�6>p���҄���3����+k@M;Z̔+��E�4��J,6NP|J������H�_dѤM:���Í!�����w�QO�z�>[��OK���i-	鳜��m�!�!���Z0�L>�O���V�	neD����[��.��zM:��H��9���9��Ri1�a��"�Q�
�s��<.���"���CX'�觟��	e���#gjٞ�+)���S�b+�!������<�ċ�b��^���񇾢M�E& �]����5�4i-P���

�W;-�4�R����㴂�S��l=�+dvÚ���\s6��!����L% 4��[z&�����tL����3�9�x�n��Ά?*�ڣ{Ժ��m�d:���Sл<+|q�v�N���r�� �w99������5`@0��	���uf��[��޾'o�g-����J���tk�Gp�� -���w��㞊za�_ T B�YQU���1�������#b!�y�PT/�F�u�X�q)�O�:ء�٫���3��}���`�;Ƞ�=&�pyt�\�0T��:Sx�d5-�BTƫ����t$��C�W;H|�wX���qWXZ�9YwC#�%-��]�6�]j%�3_�a�tN�[�k����j��Uo������,��!`=I%і������j�%���72~P���!��s������䚏��6���gW?y�u��7�δ��·{��Sg�̺�׸�%���P��!6����:�$���I��e��#@��p�N-�Ly�$Bd���5e����bY�#�>m<G'CR�m#�g��c���������㽺}�G'�w�dkm���Kܤ�U$AK�n8���"w�[+�;y�3=k��(�W-0���� �#���oe{�$�z<38?��Lm���-	��NS����U��%?=;����D�Ϲ\,3�
�-@�Cf����
VŰ�`+�3-�g����Y�=Ʊt��2I&����1�)���v���[��
U�f�g����R��UK�vӝ�@B�߉���n�u���ȷF�O����$�e2u��i�E���|lu�̥��l��.B�q�
d��	�Hň�x��f�Q�6L/@��T�?�]�K d'�����M����7�Ĭ����g��Y�/��7҇�����N����Ú�S&��*6�!c�=�Sx���k��n3g>_AZK1��l�eee��R�Dg~��U`�Xw��P(Ɂ�˪ȍ����������ְZ�����
5�ڵƜ�Yjj�$	k���7��{\'����6�Lu�T����E�4�K&��r-{��B;�u9�{b���D�b�C�)!���sYw��Rpp�)Xጕh4u~�P��i��L����';Xv������.'vv��3j)��&�\�dL�����J�o�f�t���ʌe�p�f\+C�+R.^�(�B%�U9���KĨKgf�d0?�;�d%iD5g����x��vs>����|n�����L��ӕk���̀����!C��G>�
g�#O�o���y����H��ȺEp�{PA.�Q�`3�-��������[v5H�������9Q�Z.>��z~����J_�%A�!?�>ڨ��y|w������$6"�1C�r$c�|+��z0b-g�Mo_��ᴗ�o
��v��[�C���Y�[����u�'�HxWٿ*S{�e�){������L�Z+X� ��}��UF�s���J��[(�Q8"mӪ�x�x���D�K��*��������&d+o׮ɯ0�8�R�J�따��c!�4�8}?Ai�m�R�@���|y4'%��ج�'-�����7��ܙ��T���l���r�/�Sr��6K�h���-P�L����׏�x+�e�׺h�n����ߟ��_�ش��h���Ӫ�d66S��|�h���UWu;v�`�JEN6�zen?�>2�gP;��GI���j���X*1�\�w)�^���zJ�<m�;*�>�΃��!��j���St�L{x�LZ��i!�Al����x��	�r"��I9�D��^�V��O�r�)��5��e�c'���W�p,�WUcF�=� c@�	m9�`*�'��4����=���y��;�c8�[�;	p@ۇf�=���@�'���jԼ\�8�l����椯�F4�Xi��H[��2D���ɶ!m��W���2P�B�Ѷ�17v�����6orԵo®L,O�l|lTS��W���R^�~튁��bB�~�3U[$Q^���+Dw�!���P�)�nr�}�bJ��[y"wʵ_˫ ��&��uJ�i��h6񻑤�I2#=]���f����X�z[���h	i�s}�.������9��]΍���_���4^f�)���]��ݲ�azx�%����#��Tb�;x�ǜ�.�՞��<lc=�?9�9�$�Ͻ 5Gn;���ɭd�>aN+�Xf̼����x�"M�Vq3i�GRN�h�rg0��2Xs3N�-��A[H�M�e�Z�S��/Euh���H r��Q�ﱌ�ҺG���]���SXe>řU�;����9J���L ���Bg�+��c�9KwGtӍ�>��?�e2�2�"�@��L��]2F���3�|aO�r��$���T�N�C|�/Q�K�����E+�0�C[9�W�*1K/����匿A�B8�~v=���K��B=�r�����*l�"�K�3Y1�^A,��?�y�9��p������.ƅ�ac�-�|DmN}�8]�X:������q{�)x�v����v�ID��jh����!uO "ge�_�X!+�V)��a���㏺
��%��&��/��m���i�j�|�<�cFl^��cr4�vJ`��8�Kz�`�B1��׮54�[�� `��E���?�'������=��F)ͤhf8A*\u�jq�WR�˜;pȂI���Ս�BA�x<�N1�P!I�km��*M�6��D�8)e��U����K̂������~�vV�����:�4�\-���_��J�v�Y.�Spk���Yh��:~ퟠ��9���%x]�\o~W�	̊gW^��b���x���`T9���R~�q�W��)���Xx/���u7Gu�RP1��ؑ� �`�aG�������=Е5�Ѥ�	�'�=���v����d��߮Z�x��\�G��f�L�����֫ޯR�&�ʫ�M�`a�� �@��/���^��f��iv풽N�c�0G�U\�h�&����S%�G�`�M@���j�-oa�-�I$'7���ml�� 4��ɋD�w�`�׎�O������n�C
��~�,�WE�[;j~�d�۟\�r�ؚ�O(5�!���)��|dɇyti�V� �$f�p��
� Ɖ�WF�2V�L�����9֖tw����u�=���JK_� %��F�'�WF'�i�ǂ�/�$G"�N��ڝC9hAe���=A�/znQj{鷯T��$P}���Q��]���v�Gȫ��������0~�����.?�F&�v��
������ÞE�aM⋌}��@�җc��sW�h$h2Vn���g��ɇe�p@:_@�IV�]ܚ֩�<�TX���Zg�l��xU�7�-�����:��H�m��u�U��^	o�����^�D�dT��<Lt��_�8����͆�mKb/da~�@WA��[S7�N����J�x���#h����=��i?�~�@��m�]᫝��ߕ�<�,�����o��t_�k����$@��f�в2�0G��~���^�xnH�k�`���K��vO��rk&P��2��s��[�	+)u���c�"2Y�����.c�Õ��٩u���2�*(gj-��������O���cf��T��wN9i1���ŵ�Q���eH�^u��P�\>�z��!�><���R<$��M�vu�0R��Nt+Tp�v!���)��+2$m^;4J{�c�j3�C���j��Ĥ%p�)�;*��*n&����pOԮ6��lA�������=����ncG�E�٢G\�9[!!Æ��G/���N��<~,W��E�fșjqp��D1�u�������g���*˺ć�-��Mf����?	r���B��g�K�ea���1�Ty#�e�����_��o.�|�8��bg�(̅� �<���m�wvv�?:�ז����6��� �z2�51S���*7`�&�̼�BK���r�]��a�z��� Gm$*X�_S�zJ���6sҨ�f)F}��7/��-x��h^�+�:'����lA2��wb��ݞ�]|�M�9eß}&�u��w�G].�D��j|�4u/��y��_i�ߝ�;`ۃ�ڜ�II��zR�O�:��K^�UnT�:�������m�~�9\����$�ԕ��$"���p��Y(<[S뤓6���H�������w���yyIXwv�0X{��<2E���������jǉL	F7O%���*�Z�G��/�H��}�(���8�q�le��!�7ݣђ'�z�6 v�O�Hv�-\�����&���(�u= #�8�ࠗ�Čz�X��t{�$Q��E�[���`P_�^w}�h녕����s���҄CjF`�r���]�Mm�l�/,��9��B�iu�'�)v�7�\�+�����zqO|Su��u��B�`��L��ںك��Ml.;Nk��a�uϤe�=�~>��t5�Î�p�.�sqҥ>���<��h�����[ɂk=�R�:A9��FUņ�>$iE<��)�,_���IA^;�#��):���c��e`q�&�@j�.��'�&ar��Bi��[y�����s��+H���F��B�/�w����$t�K8g��L�����rW����۫��G���f�M�O^j����K�]o�S�_�o��ʭ����K�!�g<�E¶��Ⱦ�%�cr'��/ʯ*kE��G7���I�(#��2���l�|�Z�_VJ]�wt�V�W��T���;�LFH�<�U�(��i�z}۰�;��tir���fŽVQ}ݵ=��`QY,�g�M�W�̑Ά%�{��r@2@�r���&��6���)������؇����_Ժꍿ�b�n�b����9�H��W���W}�%��!�R7V��C���/@�������2y"�R��F�'��VŃ�t�3˟th�@����%���p�"#�b��o=��t��
K��fW��4ț��i��6Y6^#b�=p	;*:?�]�;C��]}�`mB���t�%ⳎS6l�F��%�Z*�5|�8��N�]��z�Y�o�\o������x�� ��b�U\�Z�w���3��K?���t����1d��E|�d4b�j�b�.���M2�1���8�<ha���^TU�/�
`�����#^�>ͣ8TX�*ג����K� �ێ,��/��$!Y�"I�!ʽB�Ъ���l%b�l%�Q����F)0%,����������- 13�7���|X1���^Ϯ����z���^I�=I�n�\��nU�2�~i����@@�VC�O~��&����@��0^d���w1�e�L=N-]��*?�0�ڪ7��艧c�"sT��'�a�wY�1a��^w����+��?(�G[��l%,�P��qmV���m�-��DWWך|���5�~/�՚���%9�Z���8҂��ۻĮ:K>�'Q�� ['(a�����������u��)�No���ɜ�
L�v]��ߔ���Z�K\?��@����q��U��۸�G�ѡ��.��;��rZc|��em��ж�1Q�R�O���u�؂�y�*W��Z��3�
aP�ڻbD�5����<:�_�G~;xϠ�e�ct�ϩ9�N��))��LA�mT�#��@�gW����xI�y�� ƂH9�U���}#�v6���שp��$���((�17ih8��B�E-����K_��,mVC	��
������k���.EA>�F�Kq1 wJ����\8�K3Bg��������p��|�'��j������ݣC�LGˤ��U����C�܀Yvd�����p�GO�L��y��,D%�UĊ3���쁼b����J�rL�--S��u<�t�=��m�{�v)^@�7��X�}0�z������hF"�Jkz϶��b*�N�]�X�������v���ݯ䇵j:]�b�0�L��h� �8���Id�����t��㒤6]��#���v,6������i�k�\�,}"h8��6a��d�k{�1��?t��������m���o������J��u�^YK����;���I��@2���I���>~��ΐ�*��^@�ˇ��
B Pd����Qypy*��Ip�j��6���7��t�r���Wx5�쑐}E���}@v���(XO���_�T�J[}_��Oz2h"HR@��.��>*ً� 7�Z��Z,	YK�$�2W`n���ɈJ�t�56���&I�B��]4�z����ᾭ�q�'vc��j����<7�T	+�=��^F(��s��i�p�pu��M ��w!�QC�%�{�(�ӏ5��Ǧ���%�-jĺ����~��>��J�;���=K�@^cč����I��g_�^���za	e�jwn��� �A�
�k�G�F]E�A�m��j�b��[e4��b��C�Οl���#���p(a�}g�$ ��6/���1�(mX�5��}����u�g��l�0�t��y��3Y�(o��|,`��������jqT�n�N��;�v�s�'�N#-���Q�m\͞�Im�]�ID��/�!P�{;��i�:�R3 ��������$Z-0�֯�X��Z���\�@��$z���u ;E�լ �m]M���F}bZ?LV�C=Ji�/�m�q���r�u���̈́���	*���0���
���4�?��j9�î�y�KU�2�uȗ��V,!�A��hxx[ʭ_ήqH�5�a
&q�ɇ���^������M'ܳ�}�T'�D�ԎI{&@������l/��G���a�WR�cPC���²N:�\�f�5��)e�n�\v[�ս�~�n_b}՛���W�Խ-��z-�}������`���3�"�J.m+4y惡����/`έ�@�D�
��X�B
��uԯ������)$ԅ��X�^w����#�<�I�Sꔾ��h� �B���)�.Qy"�F�Q���L�{t�ژ�G�]�I��`3stT�d�^�V�!�
�7��V��3��T�<<9
/��<LC�,��kr���'�Y��ܿ���ѕ��4B� ���,5΃@i��ūp-��bSh9�n���
�l�ԪNA�����2#9��e�M*����kX�n �2��`���nT䚽�c׸?��@&�QW�nǳ�Y��%]ʵV�=�4��ٕ\�k{�`M�o"o:x8�0y�eg�پ�2��Y��`�5/kMŒ&���B��p�?�sN!J"ꎐ��=Q���9O��]��s):�IB����\P܃67cU�E~gk��Ӛ+V�ϿdCK�+iTYl4���Aԅ�І�]:��}����+���㈆y		4��R���^�T����ǖ�d�Q-F����������3$�\��o�j-���.��\W�D%9�u�4x�n �ݰ��Rxtչ����E�� M�#L����R@d�B�r�k��5���J�2�OY�`M;#����#?!�o�x]�_��:2�@יv���ܓ�__E����v��[��E�O��2���z�܄��0\V��Mk�άap�9h�-_���c��m��F&�yl1K�XMIL���kuV� �rJ3���G�R8�YZ�m�< E�F��K}7�X|��af#�W�i��Z�Ɋ�/6� wsf���w�kP�W�Q�f��0�9��=���h�eH��Q~�%�����ǵ>�7�Ӽg-�<��BB�.G|:y{�޶���p\��P"�d��~Z�,�z��ե#E/V����s�v�M�5D��"o�N��a�;v��}����~3S�n���{�X
[�Æ}_eu����Vy���.����TH>�=��r.��t�ut��W~(bX	p���|S�u�FH/iL�/��a��-��?�E�eY��&���d֎��Y@��a�K�0��{�uF��Y�����R����2���H0]/�c���*6���	̴�������������n M�2�O3߄��Bl�2�n��k\��vp�-z�~_�>)*����)��I��[��'�߷軧x�?�y���g/���wMVA�v]2Èg*u��.����6F���3�W����+$j�mWrR�[	gpq	�F߹�O]�[м�"K~8�|�.�:c?M�]J�9-<��7�R�kZ���l����DK����s��1��佴�*��v�ϲ�8�1�ͅ�g� -���<����7�2f\�هQk�F�M֡F�U��F�S*
P�d��I�V��|�J��i返���@�ؐ+f��^#1&4%�;�ŝۛ��1@a1k�vV�G�b��݉�wGR�>F�F\h,���R,�>F 1����ja�����o����͜��0��D�&��0������6Y!j[�dP�#�sV[)��i���`�x�b�����P�Xr\�/��谖��G��3|5�_��{QONn�, �K�d�+�˶�M�)��L�7��b�S1?~��@�o	����m�ҷf] ���J�o����H|�19\x�ڜ��5_���*��IQSS[�~\���W��)��Q�������o���I��O�*��R\T����E٨\Z;	;��3q	��*��q��Xѩ��xB�x�>�sq�B��o��}��{N��+I<��#�+s ~wz;�>�����T1�~��bf������کj���ZC?���^���j�.������	��S0O���G��*��\]u]�U�MJ 36=���IK���Y��a�Sj�Ϙ@�L��	��Q��7�'���Θ�"���l�� D��(n����3RY�����l=S�%7�k���X���2L�@��X%�;"��"$l?��0d��
$V�۲��t���\�V���yTlo�%D����� ��D����m��R��!lg���lz�����}��U���>�	�9W��.����<��� P3�g������Z�a�*J�F���n�K���gq�m�aX�����T�����c���4W����j+_��I��#���x�6w彣�����W�c�m��ū��<ϰ㬨�t�\;��W����@�r*�
2������#Zؔ��[���Ԧ^B^��[�V����Wq����N}�I˛��d:)Ǭ������RD/-��6T;��p�ro�nsm$YE(@AD��ob���ͺ�`[��ؗ�& c/!0(4����f�&	,E 	)�{y�X���	3�OU}����`�V$vGtjk[�[�.�Q�s��B�MhL*��W�pr*���3�k���𯆀���;�\�y�����_f�Y�3l&@���_+d齎-H��3�2q�iA����q�]�9J�V��#�@�r�\��DjuݑV���WZ�[�b�$g��J�I���aO2��<��F�||�I#�T�Z;�x�����`�zP3Y/����1b��D��;��&�dC��9�W�<�V�󍾆ZH�w��ƨ��<I�~��,)��Ҍ�8%:[+5<�g�6�u��5_8��)::��Q� ����?D������C��m���]��s�^�^k2�@�-�i���$��x�g��CB�U@(��29�W��;�;o4q�V�m��$�y��i{�ٻ�����{s�YCm�'�5&�7�)�;6���L$6�ܑ�����d��UH��'�A�Z,���n��iF�ݖ'��|)��`�x�$*�u�?__��x�'�n��Wq`��$�(��Cxk�<�\�6�������w���O�Ņ�e�ЙyL&�>�3_��� t�.w�g(���z�-z ��>c)q�}��YL��ǏN�P����U���Ɏ�[5�5H�d����j���0F�Hw��xRb\��6`R����h�����m,���d�a���7�t�؎qCn���e��=�b˵ä 2�BU��[7�"p��g�'S��zo0}W���eI'�LS,�Zܻ����8������A��p�#�|.f�2���ñ�r��5�u9�3}�M���3�|���X��̵��n�Zv��g(ǔ�]͚K;��V{2.(��F���镵��%�0�nR���LǕ�a�H����=*�V�?9y�������?�a{r#*�:�!��'J���H�А����׌T@�y��
����ٛ�<�Y\'����-�F]�r�?i��~�?A0�/��멡�!���KW��t��d�K-�o�Ʊ���Ά��lSQ�k��n�E�I�J�BB���:|�^��=� �D��J%H�S�(�Y�*p�Hfq��`��z��{��n�Yl�MT</<|��I����5dt��ﰇu/^*B��Dnǚ��[T���p�,n�koP�
��[�Q8D�����p-�qV��vyO�}����v��E���o�
��S@a�;���[�3Ln]�p1�Y�Yt|��[�7
�����ɤXI`�w�Ĝ�#_���tb1 ����|�NU�Rp���9�qo�����O����E�D�+��!�?�ޒ|<Ϡ*�d�dm�#��!���-y�\�?ފ�F4�S���&e.������D|G�Ą�M ���S����Ы�����{d	��a
O�����	��F�Yy���@aA���k�9�m\F�KW���z�%#)����9�R�XF�^l��t�E�����Tm��d�|���@7qЭ���U2�A��u����2O.�mNտϔ9�v��U�q"֊(��Ξ��/�[� �"��ٴc�"�Ȼ��t��� 1�l�bs���/\9��kN��BH�%���.�J2�\��i�q!�4/*y���W`��]j����_��>{��pd����g�+���tC_�Em��X�W��&uAA�W���ɓwR,��R����L�R!�)cQV�| ���$�] ��T4xo粰j?�����݅3ʕ�Yǩz?����.�ru��$�=����]r�ѸGmPl�b�*�f
fN/�v*�#��m��Sx�\�p���3uL��$jkA%���ע�� ���;+�wA�V� �<�=hU!oX�EF�;�2|8���	J&�������yL�a4����wE8�N9�B�2G�@8�<�Ը���u���/�z7 � �4�Y�&��{i�b�B�|�XN�cÑ�	��^�	�g��F�tJ^�
�ѹٱ�Z����[�Q6��>2.�od�����,W�r�{�C�����t��:5OO.����_R�ޝ��x�޳<��D�S~�9��AJ㺷w#^	|�P�ՠ���<)�E�H���x�S^�2�v�b��lW/�V��rK������E�u's�d�_��eٵ\����4-����x��Q�	�һ�C�C�{�"����S�Ao�����<O�3�]o�-��w���7�r;.$2�O`W�A�-H���������-?���"�#��	W���8楙�̉{����OyQ�Rn\�����4o���5�j�b3zu����u�D�9���PEa�b�2�3C��Jjb�^7�|w�/�(S��de�$�{�^c=Pg�Q��c�ys��I� G`��\y�9����3�\g�%�^T��ܫ ��u!}� 0��37�=0���p2m�~+��n-1��KT��=�a'�FP\-�v�pZi1��pt����j����7�b���������"����x���j_��!h(]��3O�D�F�O��f������{7;(8�w���ȍ�����'� ����Fr�&�H�����#��k�=2��rb3�����|���G������]:f��0Z�)�-ve�2��*Y�ŐCѾt���b��f.�/rk��}lN�]�Ȱ�l�˻�2I�wi��z&c :x�H2eW^x�+���p���.���.�_K��������ۋ0��|��}��
��u���>�)1����/�QO��@w*�Aު����Fd~7BV�4�گ����*=�6�Ƹ"^x��ǻ2w{���{���r/���m�W�9��ӎ�[�G�Ӭ�Po5 �����Q^;,�<�;�7#j�$�#�Ck���L��r��[F� ��Q��.��z������j# ����� ��DRnw�k'N�F �'�UA��.>���.Øn��eo^�ɓi`Fm��?�o�Hw��&� ��~��y���:8�V|N
�d�ȯӲao����}�&e�Q���]!�5@�[@Ω��"��b%���}K��Y>��˿�`�[�2�9�2Yh�I�W�"�Dޓ_%�5(y�<�޿�"���k���H���j�0��e�V�[q�&�ʣ���k��T�JL����q���X���gUd6�uGj@�W�{�0穡-�������t�Ɲ���ُb�p�֤tDѼ�},�J��nT�6��Y˂�<=D����ً�4�"`��a>�ǔ�T䢀v��ϼ���6���FQC�o ��_�L�<����F,���O����) �y��y[ R���C�=��[���W8=�VE����W�5�vac *e!�� ����n&��c�0T�{���ݠ"  9z��c�t���=����}�|�����\��+@��}�	�،�� ������9�V��������/,��i
/-9�̚�������sMhL��QR?i�2"���<�e��>���;�/�VH��,E�U�c^�ΫA�.��W��O��ԩg�F[�{[�xVh�`Y�>
�]�����%��GXk�]�2�//�~{�S
	�{]$x�e�X�|��y���^��!����oa��˹�	�^�?e��5ݰ5x��|���ʹ#WS�\jU�p�i�"�=�"⺎v�`Q�N|0/u�ad�}j���/�l�~�HBm�bu��n��&� ����lo�� r�+�	��w�_\��IS�e�z>�A�֖ B_$P[ڠ ��@�6J��|uc����?�5X?���X!�$��˚I�l��AM���k�)3y_�#l��{[v׸;Ao3f��;;��ٶ��|�^IPs1�\͓�H��k\�Z�cU���[��!��4��lqB�_�� ��P������;��Ϸ�j���ګ6_���[�_�(g���A[�vKVl��Nz��g(�릋Lm���%����bD�I����g=YsL#�\�,�l=ȱ����J������6�9��ܣ,������sq�r &`� ��4+��\ӳ�F�q2��U��m\���B�۟?��r~�dKW�jBb�Qj��򃶻��tr�I�WT@@JL�|>ب?\#�{�X��6? n�F�$��f;��� ��������d�����=�{�#OWv4��D	"���γ��nG� à�6��o��3���=F�$3��\��[/��	_�U:��Ơ`���G��9K۔'a���#=�=xA���j�eJ��~� :���&��+�=�����'�W"��Y����Qx��Vٗ�<�o@�rO���@��$`����c��L������v,f�o�>���":�}y@��m�����癁m!4nD�je�4�O<�����PN����e��B5�z?!�d,TSdwHNV���pF�Q�{���t���u9��a;΃:���X��RR]S�\��A �?{u��2��{�������\e���wx)���:��5��HH�xC}U<W⻗#˶; ��[|,�����9ZȔH�r���������X;0����R���7��;��9�e$d��>��ޡ����o�c9���& XP?G��9�H��bqt���3=/�2�[N�3.G��Cl�w4O��8���"G�5^�]<[�#���9����֤`�a�/�����t���彔��°u���ް��(,����鬵���1�7�3�j��,��~δ�:��R˕r�(��J���\�ǈ��v3��/K��a����FN�w�χ��:�{-L������!f�srC�֪�ߕZ	Tگ��7�O���~�Ё
n�Л����� ����?KI���1S0l.Lt=@��Y�� �QF�?]��E㺦��n����t�v�nxn'�-�y������"�|���w^;�GGof�g�f��3�Ys�ٹvv���l���dL�d@��5�aIپb�_m�wg�`:i[�}� h���Yv�5����zx���Y ��l�Pf䦦���ݥ�Rx����{���s��sn�}��rc��yO���}�hs�S�E���%W�ўOv	�H��,�4����{{9�X�{)/G�g9����amQ�иe�{�Æ����Ꮃ�v�ߏU�D9�J�^�Hdl��B�8��ˀ@$k������b��5]a������O(���q�T	�i�vLIiI��T	s�T_;�
��~�|e;K~�!$��d���s�������s��.��y.���zAe�M7�=T՛�O��~�����
w�f���ɨ{^3R2�+��
+�	��I	"JZP����9��rg���2����mN��3JՋ/�n�g���5��GT�0}�п\&�"��8׈	�;�E8�f�Oq;��^���
A\��]pq���^c��σ	��/�̖���Om��2u>�oT�_���v� ���)]�p���nn>M['�� !��!+�l^��ъy#�~Y~��gw(j��8
��I����!f?$���\aÏ�*�ru
�vvV*щ��Q���0PPK��CʭO��P���K�w�Ú�� ��-�Z��G>j���	�)+�������Cju:�	��aA"�l7�^Z*"���V��w',c���b���_�:�������U��n���˻��N�k'h|/�G�\�F�"�2��!9��O����*"\;�'��eh��ؚ�GE�X���W��r��;�VW�UlUZbt�dEbQ9n����{��R>�_�
�#ٱ��'�	��؆_��gpG�ǯG��'G��:j��cj���4R���I��'c�J �K�>��Mٝ���j��y�I�e�7o�b%�K+r��.�n�4���9̘~����иE<�[��ą?��Bs>;�A���(�#��ݧ��!O�����-@g�d�Bn����4��H�;-]�{�������=��� Λ��E�F�8�aOާŰ����v��#�ꗃ��]Zc�:�k4�P�a�Ms����VC�����S*'+g������x�b_�l��������pFP�]/	:d�-x�F>g��!E������1A(/��Ѡ���#�L��A6�թ���ڼρ��wD�S�� Wԍ)Vf�Pܢ*��[��v�R3���������6u�#�V:�o?��P@�j��!��j�՟�5�7	�ڴL���<�!J.r&���|\�y�	�'g�vhu�R,��K��g�kN������J��J�d�Y�.��/��;z�w`t�b���R��`�P�E
�]l��9�Ӂq탮�,����*!�'�� �O������!�C�Y��(�m���q�����	��"f�_��L
d�Ch�����g{�oVV��"�0��z!����i��;5������&r�զy�OTy�d��b'zuc8�:�<Rc�F�A�A�j�4~����9*��[��VH�N#L��j(�MӽM��K�rm�Ӏ�Ms=��|��DF�)&�"��ϕi�6
6�E`
f��[��R/�D�մ2DI��ߪ�db�������;6�ލw���.vdaS:d�P+|	��YɃF��R�cO�4��9&)��4)��v����7�	?7�JR���>PNy�O1�[�^nog�ɷ��t%� $}n;��{��(\B�҈n��8`Y=1�۟㝡Wa�MO5_����]��2Z�w�������`��\�Ʊ�鐑�a�i�J��0���$��N~t��g>"��~�����T1a�h��}\�4�S�>�������3r�m��*�OA&_�iq>x!g���%Q/�u�ؔ�Cx��a%�����ira�2.YAS^�U�l�?���V[�'�~|����F�C�����,մ�U�W�7s��>���{Mi��5Z�:�=}��m�0���莙��ߊ�Y�e�6D���әq���ݩ]A1�e��i�e����&=��lmn�5�KU�3.��8O�2�' cU'����oU?l�G9��!��Y�D/Rs�ot�N�y��۟���^�6��L&ߨ�֋���YG���ˀ+�{��9ޅ����O���,�|D!����˥�^�~�Qn�)*��\�CY�8O�/\ԃ)K2 �����1_�R����g���7�����\��M�vZ�JJ��j߷��
������x�@�W�٢G�����*��{h5#%�fͫ���&!���;�0��{��T���F�Jځ��qp�ßc�&M[�k�Ӎ�0Cvy*�I&&�u�_�m�'�ήW����������buJ�}�D�Vݶ+9�A�En@��y�:]T��DXE̻�RFj:!Xt�4����z��|aGC�������
w*��t�N����$���ɜ��f̶��� �O�j�-����rSE��oc|`�9[� �?���v�*�Ѳ݁�6���Z"x%����߳ T����"_���|��9L��a_i�e�Z�&e�aXUq�8[�p�����M�z�-Q�䔪g�go���j`�Q4����������oh��t���w�Fv0�����3���tHu�)�$]��"�\�m{�Ź^_='F��R}(�A��et�J^��)��oW꿘4)�@��q6G�[��ʮ�&�	���o*;m�V،%�^�iB�o��y)�1@l]v |'8��gs�����{�;5e���ea�!$��Tb�t�b?aF��W3�V�]D$���R2f��x�Ú�ml���������>�T"2.�����Hc�$D����}��
�z���l�k�@%�����a�,3���D/�x�|=D���&nڋi�:6Ǧt�Ҋ?[-j����ۖb�'�2���	�]塳;��}�;��:'�k�L��!�[�
��$��>�?�_�=�ٌ�;����ML,>�����1�|�W^�KN�	��+��e�
�E/�̀$�3$�*�y��׋��9ާI�g߸:���������r=2�a�oe'm�g$�t]C/Ul�h��48/��T�>����d���$�(�y�yvQk~ş=��2A���v c��?��?�j�O �:Z�ތ�:	�s4�Fl��q�����G�>*��Ns���7�v\څƵ++h��J;�'��wΆil�_I�O{e�MĊ�Kr�6�����#���^L��g�&���,e_��b�%o&F{9�z��O��+�a̰�q�}�r	�������~��/)\˒���ɞ�Ϛya�n����񭰍m��}��)\����%�&����a��g�w|��\�)�L���;w���z��|Ϻ����n@�ȺՏ�fvzҳX����V�CI��=Z̠��)Si�$�W	C�ɿ�?`�ۘ��.s({ob ���c����E�����m���w0��@�;�@k�x$ָ"�Xa�i�R,ee<0>��%�l|�yw
B�s�Z�=|���W�Pۉ��Y��ɿ�3L����3ū��N������vP���'����6�kT���uYeM��O�K_�ޕVn@>�z�uMc�)V�38_�N��t�Y�.F�p1��
#kbފ���{�-����x���>vw�H� $���QU�T4��>�����x^-���?&／nЭ�� ��&6j����S���\�������d�<�F~������4��e�����9��ƐC�奴�]�AJ�|��nۑ*��}�_�S�K�X0oYV%�35���&lJ8\�J�݁�w}Ao��
L�� ]����u�fx�o�P☺�����j��44�@ڕ4٧ݩ"�3૦8F˧>��E�|��� \��V����+�*5\mٸ�o�fg�`R�}}���B*0���+�O��n�pN��e��rb@��u����KgT�} �o􎊀Y�E�l���es���I��)]6�P�PY6�SxS���L��Л�����o~�x1��O<@�{��ߥ���"}1LJhB����"z�#�c� 
�{�|�e��uh��e\�FA��O,�n�=�?��ܵ阬!_�mtn$��.�QDuX��B�j+�o�{O�Ǚh�V���(�V��b�b��K�p&�J�5g�
��(.Gϝ�,�]e�� \�v"N��[g\כq��G���2�
��+�U�o�b�����ة�a��S���Gϓ�ZA�K}B�A�lw��Lp{k" ��@ᭆ�I��f��C�
H���ˠ��'ֆ����IܶwIF�@V�����6<c��7:�������(�������:����Gg�Oܓ/��ɶ��cb�h|��x�>r����Փb��+e�P����#�d�i��=?�s�(�v��]������o������h����W�z�t��P�`Q_�����/�޼�#�wl��*���5N��f*�RA���c��\Yo�3U�q��U�(hY����յ]z���1�
���&�+��ԃ�#"}�i���Wl۾u�s���[t�{�5�8W���)7����J����΄kjǩ�%R����Zi���j�%*��f��y��?)�n��:)=�]�>e䤫��.�N���1V�=�x�t�i�2�)�S4�04x�hԾ��`?�XoNG-�Tݍ)�����V���ՊnC�#�V��ķܼEk
�0��q����xF�U&�H���N��u [f��zK_G�Z�ڮy�zEd0#U�Z֠�K�oe	�f��lr�����9��@�;�k���1qL{��FL���������g���#.�Y��2������g# p )�&U�ht�t�ns� ���wِ�+�٧�o�j��!)�l���G�F�>��o[�+RQQɔ�hj���hw�Ym@t������޺g�}���qZ��
N��7b��O�Z�������,�FXW:J6�AB'�{���j�@p��}�U7_�.�U���Y��^�p~��5����`�#�nm^�J�\�\�^K�B�zs(�����w��K���yJ��>=��ʅ����
:��m���N��:o��Iz�"B�b\.{,٪7ҽ��w�\�	���5����tQ�Ȫ̬�+M��0\�'�TE��[��M�-��~R����9�2V��$�\w�nq���q�v>�����y˪zz��K_�]�g��'S�̶�M�NJ�3��4� �ͪ�OR�Tͬ�����L�Y�W�a�e�M��֔W������Z$���
�
����O�/b�]��\����77�JL|�\q(y�Q���K���t�V�6�Ě,L�{���T�M��M;���.�	qsJ�"��O�9���^�|D���oט��<c�|��t܍�I��8>�h�U�U����uLl7��ѓ��3i��E�C@�qC��7y%TнmO�f|�}��K���lƮ�	��DDQS�&� 
����v�R�5�~���)�bu�������T���'?���9��~�#��į��/}f�@:�-did�[8�.!����]G����߱(����Ր�(�>�I������EO�h�lI+�fz�T��K�V�?}j�ZJ�� ��{E�b��ӈ]L�����ֱ݈3w��N�u���h���V�,	�H�b˼�-d�gHe%�l%�)ò׈���������E��L�cJW��U��K
s�tlygggtor�?��XNDAl����F'���_���|�A-c�c�;T�k�p��J057'0��מ^�����qF4�n����Z�gx��,�ƲQ�bSvH�r	/o2~-��t��%�>dӹ��i�����^�b1��*�v���VӔx�\���d Ӂ�������$�'lm}c��saIT9DL�	h�*�77�#q�����r��-GS�����N�z�n����3�����1�v�E�G�sU������(����w�5G���{o�����^{X�ܷ`�MOΩ���$ w�Nx��wI�egI�T白�+	�P���u��<ʋ�x�1���VV,b�r��wtX��0<��G������^_S�af)��Y�<�����E_`^��J��6@��v�k4��,�F^���n���� �?��mCEA�2�N45Vc]�%���N�Q�*&3K��?3��������>��1�(}���n*�6*�c!����t�\e��k���D��^2����=Y�t���"�oRVO�CB�p�����l�����*�V9���^Ot�̪Kq��7C[�OF�D)˳��*:�E���cRߘ�
+ɝ���>�hxN�Io�?�L�p��'�硂X��N ����T~o�s��&��ț���)M^kȰd�i��W������ޯ��W&�X�yi�sy)L�.a�Y�պ�;m|'p5��"*G��4�޴-"�K�q"�����a����W�X�SU)F���������(Ժ�u�@��6�/�$yZ��_J=|1M�qp��Ūz�����^-G]���8A���V(�� /Y���*��N�����ʲ�Z�_Q�1��"w������E-��ŲgW�A4a�ّ�se"���[cK!.��m��Uv�~�eֶӮ׈-ߣn<_�Ԋ�}�w�&�Z��ƘVޞǜ�l�n��l��.�H$���|Ԍ��6q_h����g��Ɲc:
+���\�aE�Sxfu�����w��i��Y����3dy��@ ��ly�n^��ai"#�6��}����N�d��!]2i:�ĭ*�ng��醇�:N�,igrfr,���u?oʹ�������=�85m��P����o,hZ^Ӵ@ӫ<��4����=�`���_�Ϧ������O��1Ѯ�꾘ir�����\��O����ߖu֨����i����_}�3تbFg�ɏ���/2ɨ�� �C7����xiz���o�3���[����Y�6����Uq��)�U /0;4��m�O/�..�L��b�6
>R
f�}1M����q�=FHsj��'Dt�͛A��`�3��������z���9���H�C���)�� (�6�B���m��ھ4R9~�M�ylO�h�6���4lh��ms)��Tm�z�I�$�}�G�0������A�Ұ�br�I�4�/�wvj�5Zxly��?�=n�E�Qj�8��~�g&%�8���SOI����,j�/��Դ�M�k��h���t6r	{��?T/�կ�/k(i�V|4�t���qx���4���a��X�/[�ko�
����C݊���!�����x8����A?�{�y��y�� ���^�G��d6T|�f��c�����pt��;���j�07'��C���٢i�Į�Wv��QC�٪	�c�W�͉i���I!�}e2�{+�EL���B<Z�j�e��]L�^�,��zw�:ܽk�cZ�%�핮-'������[�h�n�SuCnB�o�j>֑s����،�Rv[U�����>�V�b��-/,y�?Ø�z��f羥a^�rÙM;�/5��W�Ж�	<�>f-9a�~v.��&,�Es� W��1�������x< ��&�)F�P����i�*N"���p��<�\BB�n��p �ԮaM��w�cf��&���4���=>��?O�V�T)��A� ����;@�DN1�kF��Ʉ��$���� 6 /vH��G�V�;�����s�;g]Q����L��w]� kW	�Q�D4& ���`]�Ԗ��=��t;��έ�y_�~�ݺ��c���c_���hY0�K�"���H�Elʝu�c��z���#}b:+H�/C�?��a�r}W	��>U��݄�jS����|�"�~��|�?t�{��E�����q��u��t��|fUZ�Tσ��u~'����^ x��\�@2K�������+ ������n�8>�|�dP��:��f9ejX�

Sܭ�U(�j���͛�Q��G��M����&�#��.��]5���['��$,�_�a�I�F$�����۫�c�XWM���Y�j�1��"��K�.�^���@X�߽�C/27��kc9�l:��e�s��(��P3���{�}��٣���g?Q�
'U��1�m��\�{6�ҕ7�=P��:�N�51ǪX:O���Ku���%Y�츍\ ,�:r��5H�iJ`\_z;\ޫ�H(+����s&I
y�(����q��{��r���SS<�K��TS���?c]�ö�zWPLW��B�x�J���8�$vs�}=q\�1ӛ��g։��m�5�.r?d(���}���x�/^�ԕ,�.{��_���b`�q�����a�J��8A�����mk�`���7Uɋ�a �Ș��a��l9�=w~ϙI_�#�I6���뭬j�"5���z�5Z��ZWY�@�d �Ķ���7ih�%�"2H�#`����C@�9�=�nm��v�4�F'��̙[|��>vB�xM�f��&
�t�<1>�rHl���Ŝ�������m��FgKp�~�"Zm��{�l�-v�e�}��/%���n�H�s�I�~HuR=��ӷi>@g�^As�^*��	*ϟ���	b8��/�fVw<�e��=�b��z �����ķE@ߟ�**n�e�ZNLVҿX�ݷ� r{ ة���H%��씌0�^���E�����У�%׿�Wڰ�:-���l�����Y����h
�4r_N����ϛ[����ʋ#�;Х���<�F�.�ܜ�OM�]E��[���}y��TP����Ĳ�9�K�_	="R5ap���R��&���y�qi��Y��n/��F��у�s��G0��Dye�e�[��TMqd[���V���+��D<-@\��(��Id�&N��.�B��j��]ʚ����-cs=��Mn�i[?�o�Mȷ۱2a�\y������rJ�^���3���m��AQ["򗂧��?��A�T�T���{�S�0�Ŋժ�w�啠X�Wv�Q�wZ�r�Ne-�b0���!W�����?;}lmfc15��o����Lѯ6�"���`<��VT]��L}M��T*���4�w�_~������.��Cֽ���1�R�nndU�G�0�1'�i.x�Y�*��~._�hW=��.�=�P�ˢ�;���E��8ܑx�A6�V А�	��{x��4����>g4�	�]\.-�\{��Dɭ�
�=�D�;N(��ڞ���B=��+5�����ީ�_��*b���iG��Wl���D�z-2�d�>`H�$�#!)�!4vQQ����������oܘu0�p��B'�4���4+U��w?X��6�����|g~�|�����g	����w��kI�(��q��i%�b���D��q��O5�U�%��0%��Xqu���-زq�61����O5-�fi����k��'�P��g'�ce�׃.�S;eI3�MO�f�g�����n�i����p�SRmj%O-G4�������Zhc{�>j0���D��e�rѦ�v��9��Dp��
Mo��yO�WF��#6�j(Six[�����M��׼��$� �*{�UPI�l�@_lw��[�5\BD�8�A��h�֐@;un�~�.�C ��@(!.	�	E�.v��e.64W���.QQ�-��\�0�O�Ą��|��Y�gFS�4���d_>��	�E���v�D���N�q�?k��ɱ��K�]O&6������D���<
�L�٣��.[�������c~À}U$���e�C��#�z�j�)�M� �6��~	|���'l}2^%v�zRҮ��Y��?9�#z�7^�P#r�J��ޯ_��:���s��?
�X�'�j�Z;`9����+���Tl�m��Nf�����ax��K���>��1�n�)���L�A-/���,��l��, Jf�z��{�"���jTe���fKZ�~��q�2�_i���R��}�4�'����"PPX}�O*4��x���T���H���DnF���~'n�B���A���� F�e����C�	Ա�6���
�~>���rF�٧P'Hמh�qs��W1*����[�������w�0�}N؟�C�|{ҥ�ŏ�[Y�[���gz%U�꥘��z�$�T�f�:�ɗF%8�cVɔ���`y��ٱG�[�{CkUش��'���ɟ{�1'��mJ1��9aͪ��B�Ͱ�"M��zI��4�Ų�v5�+}>�`X��d��M���8W^49b�Ӫ���p��Z����U��ۣ�5�Ϋ~��g{$����'s�S��
�r�ʵ����1��})�K�K���Ʈ �Q�ROX$��ʿgC6��ٶ��i�3�l��O��7���=X0jQ_Ѡ�����MUx6�����|���X&^H́7�
�L��D�Mr���V[�QX��
b7�5.df�kU����M�S?�X�'�G�t旲J���gR�3�>WO1�Q�szȘ��u��-�J?�ke�)��?ԗé�?3:��IIQYNwH�H����������������U#�5�K���]h>���#<i�Y�"�S�d�5�,����7:��AF��ӓ�^�����p�m���fYj���Kϣ�+�C5>��jW��պb%��/EOic�.�R�B[A5���3���
3b����ձgKB��r!G�����<u���.�]I���W���jE�k�._X�`�3�H���IL�B��b.��*�B��A�O1ș��~�vc��p�̏�-l�$�Ke�e_�jR�#Y��\l槬H�4�צ|�#��[#5��Q������4�&��(f-�\d;WੌY�Q�Q<n��Mml�+)���p��u�|h�[٫A�x�@��DٿX2''��ӓ�f2���_N-��`㕟��*��[,���=9h��C��J���F��:P0�M�����������`�@B�S��@}ųFܗ@�JX��o����%T�%
�8nI����.�J�9O���&��cփ[�;g��\�7�au�����&kb��U�����`���D�&�P|�NL��Р��C,���e]�*���.�5[������v
���}���lmR�͛vR�X�"V���u�;�IB��/%<���.�_O�(
w=�LyU���Ù�\<W[�1�	���&���#�&E���ĉ���N�s2��-�1Q�`�Y� ����pi�V�G
�z����r�mte;��вԍ@���V��SUwᏦn+��s�{q$w~�o
���u��A2��֧��Y�^Н��)�"W�6M���W3�X�u�i`����Ŕ�%�����\qlX��P���YhFV[:�s4��.� o�nv'��iy'�8��Np����ɧ�<�����<� ���w#$Ď���D�y��+�+�["�8<�>b*ğ��UΜϟ��(���2
��i���bwr
�m`���c�}�2��
2����@銕:m��C,�g3�{{u�����q,1t������I��"�h7��̺���_Q*��6��c*g�oȵ��i�(�V���۵�A�gx<K|����ܶq����N�������\�ӭ��W~P���2b�A�Щ���b��ѷ�&��(�Ri���5j'뻝�����JT�z#�, ����;
��p4Փ�r�|5�7� ")�C��K�H�PNt�l슦�z�
hB�����o
Ym ��V��]�^�x��_��l��&�x&E�l�j�$����{��k��G���z��������%�\&�T����;j���������?6����fRN�Q��S1G�1oq"�ĲX;	a��_(2�Vd�<ۍ�Ze�?A�}�\7�}��lH�iG����QD��X�yFG�K�ǀB ��BЗ�����S���h�WK�_t �C��!���G�E��ޖJ�O��o{�������z^�Kc�4"KfI����������H!��b�m��ub@�jh�&��Y�ڕ���-�����{�޸�]{$�H�@��`<�
��T��͌|ۘ�}�i������]�q�R��p������F��\C�����LB�ȚܔZ"�B�#�ƃ^�Iܨ*/��SE���r$g��f�M��F�mMD0y9��$�݁�OJw�� �#���*��.������
�՚5d�;w�I�7| ���`qj�$�܌q[�%��Bt�?��*,�"a<��^����5g������<�ug%r]
����Ҧ���z�l�nl���Z�Ը35���Xl�����[.i왙�f3�� ��˾9u���>(3���1�ٍT(Tء�T�s���oSB�~�ӊ����Ѥ]��΍�=,//���3+�F3��9o6-���w�{�����]/��K2�����܇L�7�A	�x��I�K%ץ�1\]�D�H�&-��*����O0+nl�"4����1f"2ۦ׳3˵������M����[ٯ[���_�+����]}�B�y��!x�c :����
6���-9��aY<GR!*2��q���e�E��Vc�Q^9�?B��w�4��mȥ���!�tu�<�U�[��Wײ�_]Ӆn#x���0:Kã�r��i���[��+��癔�0�=HUs�E�	QP�ӹ��E(���^d��D�iU����k�{�� {�?i�|ÊP���a��yZa��4)�#m2˱��ƉMk.���־�Z�<N�{LꞱ/��,/����X]�[�,��/�6`���'C�|al�_��=������D���@;��C��i�!´s���t@�����mJJ.�׼�bz%^�YNg�t�����9#H��G��(�)��(y�S�ӿ;o�yQ�[ Kba�*�8���5�����\����O�3,�kP�-F���1v����ܕ��4��K�=����$���iNK����+%v���n4���+۔䜄������f�{~��J�!I>��d�=�M��'�^�e�yx�Nu����<���1�_C�����}��956**�����~{g���v�m�¨��Ն`��ZO���ىD"������
~Mq�n�q޳�o�`
��S܂�'�->�y�%�L��_5�3�����>##C�)��R�Ѳ�>:&f4��Cِ�"�&�z���b�pggg>Hc0��ʋ/X?���6�����_i���������0��0�p%�w �v���C.����?<�������W����ꥩi���x.~��]���3���\�-����F�U��X0��^W����r]P���G.<S��ݙ(нqd�PO�K���"�"��+gv�����w1		0���D
�f��.IvEf�$��#��{�������J��ûFϟ�W^dLv�q5�QRZ*�
��Y����7��,0bk�0Le��FGg��)�0�lwr��v���.�wFrE�E�M� ��0�G��;���y[��1���+�c��+�44\��p�h�3[A��aj_�z�V���Bz��57��~�6�c�	�>55o߿�Hy��B�"���K�[\6�i/�������`'��U��E� �?�Q��ty�4W����{,R��'�ˢxg ����{���	�JJ��������V�����bӀ;�_C%����rT��#ݾY(e�؎A^ߍH�B�|
��[4���A�R^\5H����!�s�=�̔�����w3��W�.%��OY<���6LNA��u�,!�[p-���?ن�U�t�D�w|g���Or�[���ڲU�^�N+h8���hg�/��<a�ׯ�������E��[m�.�?	��A�� ��ۈ��y��?9麿!g�EWR�f�c�	X<)Ĭ-��t�h���V����rz����0�/Lth	Wwo��A1>��s�䉡�&&�������-)��0N%=�|o}�Ts��{[�H7�)����o"R꯲>���Z���Cn���y���z-�DEG�B��^}#���H�,A��Yv�;�ۤ�
ȕ�A��̕�HM��
��ͤ��O�A�
\�n7��H
����$u��K���$a0o��c���c��U/�8�c ����[��H"�ߘ.{��N�Ĝ��J�e��ћX|b�}g2��:�_�tZ����7�}r�2�C�~v7o��Y�����	��s���Ň�zol�,�Z�q}RȆ�5��W�/ffd:7t����l	���kx�Myw�N�&�w�����I�_A�\����a�V�S�߯)���%Z~kM�5��p6�6CF��ޕ���.��//+��ɑ�m���)�˫Y[#����k� ����c{w7�|HF#����BX>���A2���5'Ǉщ�}eu�
��y8� ���, �?k)(|������r����505�p��Z�b��}8$!�k��1yR ���z�� � ��^5g��V��/�eZ����' ����]]��	I�l��81lׯX5����@s�����,ׯ@|����'?܂.� ���C";���7��b�D��������A���e��6X�<������~'��g[k��ش8�r<������Vz�-O�dhg�����r�30�0Ը�?3H������}�z,��pRDꐈ
�!{S�<^��'N!�ۃ�8� #/�F��F �X桦��Pڋ/�ZZ�iоT���:��`�����ɏTփyz
rr��1����5q#�- �d9���v� �^=C�er$w�_%�ڈ҇ư�1)�,�D��n�~�l�p۬Z���E�"�+e?�̷J F̊����Qں(X�S,���g3kyy��^�_f�ANEe�h�V�^�v��h���}���5L!1��d��I]A�W��^r�* "����G���}�x �]7;�]����b���ؾ�X΁~�� ��g���Y��ׯ�h�J�D�������9���	o�a1�?�����A�o� [��E� �w�c�Q��{?���sm��/�YV������XE -Z��8�@r���l��V�ENN���Q#�|��*���ÂժirsssB�P��,V��Q+�{��\�	���l�qq)��[��9ޟ�/Ԙ��L`i_���;ޏ)dcg�R >�0�z�6� A��P�O~<ow(����U�D�0bJ�ޖ�`jH�����ףȘ�lŞ�+���2~�zlp5���	�Z�0eK�z/0f֝r���|������@�^��߼�]�_�K�H<F��nJ���纒s�P����%(� ;*���5��{����3��i�ͽ�=\����ht��v�F��|�{�,��z�������%������#KK��W%	$D��i����ז��,�s�:�mJ�����c��C��z׏(�<�����#D��Bo�<8����;Z����&�R���֎p.�W>d�KF��t >��zf�*#0��G�T$� l�~y{{d��v�oi ��5Rj���G ������c���aQ.�������(�$�$-��H���>hdYn����sT��l��dm��j'\'i 6�ع�U���ө��7i�L��3/�0����j4Nn�w����.@��0�ȩ����
�a#����˭�Z�r��O�����rG�u���iw)Rk�3,!���a <�)i]q�-�+�������r,͸ދ�g<�Iq+s$C��i4�ߟ�h_#��g��t���!��l���@�R�i�P��K@�Y:�U���Υsa)i���XB��77��}}�_~v��{��\�9gf�����ة����힄��㽒c���<}Za���+u=k^H@ ,����L�ww�u��h�=PkdL
�[5j�����0iTE"1e���CzI��� ��������)�4����;��x��h���fhm]1�Dշ%���i�1�z9kk�4������?%Zɱ��Q�6��g������x�#J��Q]�z���r'E�WLO0?)�w��Y%��2K�,HB��\�4Da0[7[ί$�DGG#7��f�w������_�Խ��b��࿷�3���	0Μ���oP'	;�U��ăΊs��Q;fq
���+����^���n��Ӝ٫歟��d�D�:[˂�X��o�����Y�P����	֮{�zc��U��� z���"�]ޞz|`N'�%��������Kos�z��kKat����q�����#��3�N���1��#ݜ��7�>{�1aL�7n�|>豴 ?��bhC�\YuJ��&9|�����m�zC	:Q��h,�ڧH@D�m'>�)5�#	\�04,�}o�-��������[�33���1s㞫b4�� FDW��}F*-kg��p(��ID����<��-3��V����{�m�Zl�#f���f�}C�v�P]G���K ���\�ǖ���3�+..U)/&	/ہ�$��4D�������\�:�#/e�m��ҷr`d�ʔ%r�F�B#hK�����Y�}�8���;�ش�2��p�Q���������A]� �p�.װ�vGeJ2���i+x�U��SZ��F�jt�Z*ae�׋��`n|o,��S��(%Y�����A$�ra�y(c�Ĕ"����}vM�����#�mm.��(C����	��Ŕ�Ə�$U�uYRJF
�5Z���=�A��w@<��
�`�<)��<ĘGg�C����V����}:[��6PSS�V�T�S���7��"��3�����mqyy�ؤ��ֲva�d�n�՞��!���e;z��ׂ�.:�+�s�I�2���eѴ�
W;�E�o���L�_~��*r,ߙ�	��]I¼�0�f��~�$R�SY�-Z���&�"x<\i�֛��0Mf��&��P�����n�9Z�
�1�@��QQdk�U^^�>�� �d�Z��8�?l���
2���]r��nn��եN
��O��G���a�_��'b��Π{s���8�P9�ta��i�DQ�E���/��y��uy$b�X��8p]eX��|`����\*&�3�ܖ�Q^M�vg,7Y�p��QA�Q�^Ȑ�_ߐ[Q	�{�0L�?$Bُ���ގ1u�ӹ�e:�7b��Ɨ������)흩}��nP�.�'���rd�b+�o'�r�"0��ZaU H��WX���D�����9p��^�^��T[�����HĔ?1�s�j�f�JW��򋺭���%��qI�h%Q���#��M��$��?�^6�j�,Q}U�9��t+Q�����$P1�ۜ;�;�Ő]}?s��O�UV����x�_���bg�m�w�#�s�����J��$���w�.\�r�֦qΛNu����(湥=&n��z����ꨞ�^�����d����Bb�O�^5�����}����{�.a�TV�cي+�����\7�'pڍ_\��N90���?�w�_翍��w&?��*��z=W�~�L�f�{YKS3a�q��'�GG�O��gp߀�/㜆��g���������9���x+�.�4)G�K&�z��b�A���$����x�4���D����7~KK֦ff�)d�$+��۶��{*


��4yUw�ڙ�$ZH�AZk�q�������.�7�#��`i�=:���q�c�]�K��W�T���ފ������,9g�w�g���y�q;��K��cȝ1�kso�؀���U��3e�c:g�f:c1Q�7�w�BF�&����������<�Tq�n���¥<����l6����jQ�B ���hhdo�����>;� l��T�Xd��m���k�hLv�d�s���W[�F�6]�����{Ƕ6sU�@�C�?��F�N�h����kL���&�O`q���{t��k>����U�5I�\��2��-p(C���Z�gנ�����ڜ``��g#��x�@3��UlհU}��Z+��ԂYt�(%��Q-+0Ԙ\Ԛ��V��㫊N���ߌ���xwN�^P�K2�����g4����C�$��5}�PhtAFƃ��׮���[���.�7���z���9���a򡆺�<��(�-o!���gYQi�SA�e\tI��q���� ��!���g�ZG���V��sS(�Ew�Ы�{��2����y���򋋻s��_�1�geee�@����J||�����Q���P���*��Ά��7J B
�C�G*0t�r�tS������ƽ<g�䟓�jM�7u���5z�����X�܊M�t�R�P����"�I����;�%(8Xع�Dw���B���X��+�184��O��*���%b\��A4�L�0�%�t63'a.����8�K%��ƿ���lsF1��(� �R���[�3ZzX�c��Lr����+η��~�9G�e&�Q%k����,a%O������տ�`���\�����}}��������,&�����Y�;��%��߾6�L�5k��5Z^X�W���@��<X��H|Τ[�{� ���J�LXWt鬝��#�Hn��{���/��8h�$	<��<7����͎��3� g(��41�趴��~j��M�2a���E���\�PA��ٮ��$�n�/��&<1}ڴ�#'Ɣ���3�tb�1�7o��<o�f������e
SM���̏~����H�������� Ԕ���1%S(,4�^ef�ۊk��A�/�x�
��q����3�����\�CSZ3��/t�z4��Z?����8��c��sk�NJ��kOGG��YYپ��Έx{A������rOr�'<�9��r�j��ovM�c����F p�!54����.p�&�?;r��?_+��$�䶓SS�=Օo�Y2��4;+��v�``�g�}�ll� ��(`������=qrZ���XQQP����R�yYY#YU���b�g^\Z�hY 3O�ɇ;�yg!�Q|�a1����m6�.9�_'��C
��걸a nL���m~�}�R�/V? $$�oH��@��#�1��������(+K>�P322�-9�|}��D���]�u�\h�^jjju���}��i�Z>�o�P�CdsP�
��|Z***$�.�3��S4�/�̸�I^~���:����ꊒ�}��g/ ��V"��ɞ����t;�KX��3��_=��^��Y�]���pxT�y
�Z�ݫ0���	C!5�������gd�;�q����M��R�r�7�&��ݫd�#Co�"����7�Q�ۍ�ʗDƯ����CWV��Y?O#��u�fkO��W����n��d>R ������Z��,�Ç�̓�
�6Nt,�ā}�:�sF=����e�,�6٪�cj�ι�=�{*f�ך�7�?AP <��V�\���9����X�%s%#�}����W�wy�Dp4觊G]�իtn��&������b���1��-��"V5�&pv��l�P���6�r�� ���9KH�;,��`�=������r��oO��yq��CMU�����6���в���%��2_9J���K����F��~�A a�2��>�I�G��G��s��B��m�V#����bn9�ua�~��&?���$��۱21	E���lk�$d�U�_:
ḣv��x���b���喳�(х.�Uh+�D�hz�o<�b�g � ���yc����[�b�2�O>��a�^__���a<�]�x��a>����|��?��&}����i���R�_7hY�1&��?�@���8^�[]A�x�����X�Evv���Oo�iv�P�Xr_{���K�+���K��Z�a�s�N1�P��;�M�3���v]�r=�}���*����3��u���߀���.]��nh�*	����}x`��]U��{�@�CUE g�e�2.K�� �~��9���4�����X��������,���c�_�����ME�"�#�A�讟S�[q?�{��㖗�V��n7T��2>�**�r,�!vvv^؍755�F311��׏�t����OӸ㔇�@�cp��s�
����*�`�0מ��>����Ci�c����H�d�RF����ş���݋�>�fn�Z�u�Gu��R/:WY���::��:�O��n������^ K�1�D����	R���R�M>޽۶žG�Լf!�er�P	;fEDD���/?��s���XvCJ�J˝�0<���jt,��o�G#2?r�jR�R�!p�_�v�@�4q���{�l�����K�]e����Zʚ�J,�0����>����0�^��1�<�	M?�>>ޛ���(q�m憬����q���w(F�ٹ�m���s],,-��J �� �!bz�D�c!۶�=��p��T�#�Hל�;�L�K�,?�L,&���A��ϟv������
ŝh+]�S+x7�U��2s's�������k�m/�C�iY*����֟�c�{1�$!Y����Yl���0��5��d�og����� �zř����W�"�P�l�ߏ���T.$��7ꗠ4Uh[;�N;����+%�tg��s^�5K/�_���DϞ�;�E��_���`H�h���Uuu�j��x��["�98������L�۠����O�C'�<�x&~�}����S ��g]�:�4CЫ�ߚ�m���+��\�u{]�������Ko(D�'�������1�!�5���TZN=�}��K�/ķ6�r�J�0��7�i�D��ت�=�������e_��7(��$�ZR�W��u���&(<�t|�z��`m�QV��_/�a�d�9#��tɋ�6��Ŷ�"�����iR<Iʌ��A��5�\�bҁ/��� ,��w��m��6����|�`=C	߾)@�K����I�\��J�^�7J��+�\�z�����Fd��S��~��/ᆊ*�~||E
�����3#qq�ٹ��qm)���O����:nW ��ӗ�A�|���{�Sx���Z�t]�
e�<�0�G�{R(��ϜI(��[���jTB�A�!O%3*&f֕Ik	[��l��/(Y�������G1yihj��s�4>���F�����5�ϥ6������Ľ�(������H̥��\ۀ�y�	��^���PJ��:7-��.æ��۰�N�
�P��XCZ�m9.��#�X0��Qm�u�d���D��PS3.��<����A���z�>���W.�JNl��J�Ґ�n��1V�&���^����������LG'���]Z�+@|-�5���FG����.q��L�u����uYwfn�s�e��#���&`~�{�ɢ�I_DDu���m$����EE.��ő�`�U������.k�G�����gDm���R���|§˶t���c~����N�ފ_�\2Ov���u�IPǘ��cs1�a�m��7���ޠ���x�Ժ�H?Ҝ�\=�ma��}�3:.΢ �3N�^\���0)�ۯ��V��Ýw�E�1�n��xxE�������GP�n��:>����)m�6�QM3�2o�b��Ś��o������af!9�����e� p�F���5$.�a�N3����c���<��ɓC��{�%���#�1�p�b��T�a��XD[��,�x��5�Jԏ�t)Z�'�'��ј�������F�PTl,�+�_qHCCc�=+[>4 �Ɏ_�b�Z��������l���|��U/ў����Ӂ61~͙��K*k}? ������|7�1�*RsOP�����m|���5��_�,�ju��8������b�a��Bn���mѨ/��=�6 ��?|�xF��^�.A�j��ՙ�vr^���X4��~u��V��7Ԝ+*�A)\�E�|��'�l�E�u�Z��*�ÿ��|^�,XD��촶�����ڱ�I�Rg��Z}Iy��}Z���\5�+Ub��D��z$ե'��ӡ�P�$��S,z�wV���By�e^�Q�N�U �lF*U���܎w���������p�=ru�˃9�4���ޛ�����8�O(���m��KM^�eJ��{�l9�m��ûq��$�z�$���zRl
��XX���n�+M�>j�v�5չ�׮\�D�5H��� �
-H�e�|��ł5d�B��6�ￂr$������ؖF�%Q����Y�0��d'�՛��N��y�{�k>sQR��1����UwO>E[i=|�N���P��I@�\o}X����7�t���J̕��C2��Z�5C��*'�O�eee"G;S�蹹9A\����!~Y:�Ҩ��ş��r�Q�~'Joi`dgr�υw汹��M������ ��?���	 �kB�6Xiܷu��a���3OOo�1�uŀKoc��w?;ڜ�i��������M>\�~��0�B�P	.��`�Ք�[,��4�@�i�(�kdh�(u�}�q���ӽ7��i��G\��C� �T}�U�][�h��4���QQ��ͭ�e�]%��k�C2�v�S�4׭!+x&�S\�@�s��ԯ�A5e�>�������Ju Q6C¢�K�»C �@Ã��x��&�&F��^�OtE�}��x�����=��?�M[厦MOf��וּ ���ck<�ا`��PYZZB��Z9e{��cwfh=G�`�����k/��,}t�?π��� ��]'���i2��.�j+���e��<�l�r1���n�Б6n�Ⱦdx�t�xҵ�BO��?�����o��\\�Um��E�/)�^�V�
XR�'GGF{./WTٍ���-y{�n1ݝg/���h֧��cvv�Nq���kp�^�cv��X�'�� �y�`�}?�V�b;k���Z':���Z�'b7�٧b�e���a�Ϊ��Μc#�����+*B�ٔt~��0�hm���B�-����CV�5ؒ���i��|�m��3{%�#�|P~P�~Go�~DDD�γ>�]3��c�z�����Ei��i#��Iė�������/č9xO'�E2����ѝb��a.�X����/M��=�;�e%5(m,�r�T�Bڧ�����܍5:8��GGG��؁YX��w��v����H���
 q���:�^�)b���,z�n�}kԚZ�ۣ����*��*�����x��nǳd6�,SJF^�j̎c|k�*[�����������O��T�(&�w���2�``(��w"lhU�E��#�ڰ9�Gt�t��g��-f�����B�m�b���&[;�X�G��mm�3^�$49 ~��C^}2#�h�o~u����әw��D�h���� `�5���>��%����W�o��eG�� g߾}�1�꼍u�$FEeA-F��!���&��< ��XCBU#.>�Z��j������p.շ��� "��>�)&�ﻏ6b���-�W�А!j���<�z�4XKĘG��RY���p�t�JS�8g�Ϟ%�d\�
�l+*�?�L������jx՟�u3k���ׅ��L�bao7��AC�Ǘ����;,d򑉷�`��}�.����@a$�+�&�@i��k�4)6�x���6�]p��U� £s�4Ź_�+����BF��!��&`7b8%�^;� �Qi�y%%���P�h`	�Y~^�c����8q�=���|9eeD�
��+�::9�簾'����!�D��Oz���,%a�ElA���jq7�go�߈�;������
��Z�R'^�����W�^�D�`G���?�H�X�/�k���,T�'���F��R�P���0o3�ۦCW}�.~(e=��D��4}��y~ԩ�%9X�4wuy���*���K/8�k�S;�M��@4z�#~|f$� xZ�xN�-�F~�n�P�S���f�ʭ�K�_%�b�Y�ؘ�8�acc���"5x;�?i��DI�(�ߌ�,9O�)gp��Q�7ܦ��m������;b�o!!iK��m��f��8`�n4���97oy���[p�n�~�O��O�/��*��}T~����e����O��&��X	1��r�~��g*�]P'��4�Q�U�_���u�6�9������z���щV�h2�Y ��A�<��_����ׯ_��g?]�V��Nv�Kv[���D��S�=��ڭ�~��A��9o��=ū��/�����C�v:�$�V��n\�u_��3p��
F�#���;-����Qv}��2ڼ�ή�E������k+����?o@Y+�B{w�2Z��po�S_&�����s���މ����vq]]���E�z�,o��a���RDD�%싩P(�h�^��#�����~��&�^�vc��~�X$'$���������L��*���J�zw��L05X�qo�b����F@�����R2�m̽}kp�o}�h	Bϟ/5<T����_m2�Y���i�ƽ�fл�6��\>��4�Е$�V�t���}C@@Ӹ-�Xt��eB������t�������`�[�5������X�Z:��.�#Z!%��!*��j(e��_��s|�4E,���̓����u�X�������'�,��P`��G�5�q]��v�p���h��Pih'@�L)�UUU���
��1@g��zr�k�	cl���c�Pgp<�9$EK��89ݰ.� p�<�JnPpp82G&�^d.ɉ�uI;;7W�cU�L,�{T����^�-~X��vZ�;*�m�c`j���X������*@������d��~�,1��旃:��G��@kUiїaV��M��E�xڪ^.~�������zΰ@�?5-�~~؍�S5~/�r��N�6@�d%��@�cq�E6��h�9+��~
���2���៉B��1<�T�#괪*��5�U�99����~�hF�8��Eѥ�����eJ�����,Y��(��^�}� ��nb@ðid��,3k���|3��_*�덙>�n:ևz7�%������5��E��~bjj꧝�PL�i5ߛ^�����G4A���*�F�.AAA�:�]�~ �#��+IJJ�:�$���q��ˣ�v	�`[ۏ �.\�k����рF�v��p��߯�{���-y}�����atR�����#��W�5�l�w�#=O)H}2D��g�n���&]L,�0_��
/�NH�䐵��T2���<�}t��O]�����;Tl��{��1e��a�:�{&V��|E�Tn�� ���#����=X�8X���2-���Й�2���U�����J�l�7�������5����j\�Z9�%��Yf ��ZC�hML����iS3��'��)B.-�_�����r
ҍ�</~ �q��g����B$w���&�����S��"�҆��8����;���*�P`D�8\�뱵D5�<�]��U��,���???�W����$�w�y�l	P��ր�Ϯ)�)",��·ՇY"��#_<	s짠͕��@/g9H���4��M$�ώ���w*{��� �>�q۱E
����c�|9p�,˨G�3;D���sY��W:+�-����UZt���L#����׹D����Ÿ��~+�S�ɾ[�wuw̯��y(?�z�©`a��q���{��$���J�A���� z��(ʶ��çO�}7�,!�Aع�~%���D�6����oC�k�B�[�h�������|�j�#R�H�D�|��!���ˌ9��\t��ِ��p��=ܿdܰ��1�72��O����"W��)%��l�5�o4�����{�9��
�Xϰ���H����-�=}�w�}�ۗ/�y4$8o�t�٥H�:�vA��)B���޶{^�	���|�AW/nDr��mQK����i,� ��)�#��i�~��ut�7����G`%��+�ak�P��y��W/9洴�pP��h����t�7��3W����%�ħStU�թф�7���*�K�kM�kb}���\�E��!�(���� ���Y��U�(dS���Ä�UZ2�s��s����[�2PH��M�vK��JD��(��ɟ;��J�kW�C�~*���1ş��EP���-�X�Y�)�C(Q�*���S����jjhd���>�`_��4ڏr|��[�=�+f�� ��������||�p����6\�j���lؤ·}���_��U+��v�mX$f頓��t�K�/S���<A{�0N#����yt&�wA�рqcw誳���r7O�v/i*6 v%~Ԙr7���
l`.���eg'�'Y�w��T��@c�W�b]��|=�>���: +G�(�|�r�3d#Y,���7$|7QP�:�����To��Xnt���q1
���1�BN��:�4��c����N��c��!�N;1��+�kK�@S�x�	����1��C�{Q����х��TŬ�<����Dj;��0�`������	�>�l�>ɖE���ܾgn;����bȟ$��>@���_��h&��J/�k���ߩ����-�E�zaº~�)����1v^�Bå��ah.��u�J�
�������(6��ł�Oo���Qq�	l��[K}@睻p�Fu��e����'a�ӈ����x�'����q�r���E�8"l�z��GJ1w�?RQGw�*���!�ZVld>�2���ph�����W�sJD����� $��"J�JZ��$\�r��w�U�e�&+Z��~��O����'�s�� ���(O���..��VL�kih�IH2xo|ߛg����ai���=O�i���`Wd�/�ǆ�KD�lOߍ�8~�4���5��O(���~��&WʘC)�{B��v�a��'ڥ@;3�C�O��w�}L�;:9o��31⩶fA�!��Q
�2K�.|�B�2Ԋ� Iu�Q�w�b�3w(7��i��R�g��ְ4S_�ؘ�iQ�P��5r�Q�^Hqڷ�sfD[��v�G1��<����m5�Q4�$!h�rp��hTu��Ǌ����*�?��M��x~q��l�g�Ib�?Eبs{���{l���t���ԛFC�@�K~������`Iw�<=DZ��|�^�������0
�V����E\�jjj̖��7o�a�j,X!cjk�8���E1>PR���t�$Z���w�Ξ���	XO
W�C�����-���%��Wd����m�^����Uz�4�hE�̩I������f��j �B�딠�7��x���#m=�ͦ�k�����!�]
����	�u$og<��Żt����G��b�����'���T����|{�3�e5����B�T�e]�8v4[���~�����"k�Ey�v5��z�i�x9����zš�JG�Jp�V6h�Z.l�L�3-T%����@�طT�������$oW���>UŊ+��-�*����܂��h�͛T9Y�+��Y��t,ߙ�'������|uF��v�m������rB�@�ʊ��dfa���RQ�1��2��"�������g^` ,q��$�]���������eeT�Р�p-�5A�i4
5��e��Z��o�3�j�J'}� Lɲk$�>HQQ=�����+k2�����V�^���D~�f'�cf�H�[�N���m�y��L���j�ԻV�E�G2-nw�n�`M���M���E�d���
�(�dLц�'���J.���6t�^��c�VЩ�J��4y[A���6^������I��z�$�W���`(ȫJ�R��^���B���F��c�ys�o��Jg?F*��0��?�~��N��C����w���F���F�N�ɢUNsJ��7ђ��&'�_�v���dgԏ�7��f��O0��u/:Oayй�����G�Mv|w��Vl4y���]ZY3�`1����{���u�2�[C����t�����%���<�=�OD�0-���Z��n���&m�m��"y?�G��O�xގ��b�7z�S�k��'>����ȝ;SL]���n��t�����1�5������f�+�FX��^���q��ѧ�0A�q݁X��p���`���*ѬH%1��f���R��y@�a��ٗي��欟��o�x�&�Œ���k�iД���0�@�P)/�qt:�4��!��ɯ?����-g��!<�C��Ŭi�#}�3g�P�r����*{��%��1�9y#ݷ<�s���C:"��$��Iņ<s�DWZ�w�\6�7j�Q�E�&M�5\"_O��Ú�dC���_����:�܇�[+�S��]�Ll/�$��39njj�%�7}���K�Po��__�<��2���{���}X�+k���n���*Ņ�p7���bu��M�mV.��,����u/{�㥊�B�ѓ#2e�
Lp]�_�)��>�k�*��縇�8nc�<Ǥ�n7�>����H� 5��mf�f�]S���=�>dc�����Wm��
��#G�d��ͷ]�PM�i�3+�N�O��W��8�Ǟ�#���=�~O�[ߟ_�<j]�=�z�����-�Dad�VƊo�W�l^�g�?�ua/��(_�hƳ�Y��Wb�FNn,���m����Fj��0�x��虧/W�xļR�qC����h��������8l�8�T������c^%I��s��c������.��K�q���ϫ���+A>�="���$�%�r���]�1߲��)�L����1���ҭ�Q�y^(hb����r��q_�q�|J��b��W\{Q�(>~�"�:܇2�.y%l)��,*_�[	<��AH�����ҕh��������Xw�<Y\�KI��#���=�9��g�V�_�y	Z+��e������Lr�'G�Ep�y�-^F)֫]ۇ��jY���va�ha�8���5t�����94��.|Ѿjfa�nCl1��8T�6 ��P�L�k�:n˭PqL)ds�ՐT�0V�2t~Hǉ��0mwu�S^z�|wF+֢���K���3T�z�D�1�%;<���$��pM��D��(�UFX�-G{�b�V���%�7���j�bX0�`Qn�l@����i�24�(�*���W�|�A�b�v��˫v���������qNξ�P���Vt�������]km]�n��Q�bIM���s{Ɓ�CA�6��B�G��Ӑ�����Wi�N�q&'��S~�s�2��w6��3��N؝6�+Z�:���oc��E-��Z)���4�E@�
�0Vߪ�5�Z�-�S���
=x;l����K[ ^�r���{��.qD���D��k��X��uU�3�bH5A tޕ7�w��¦#pʫW-�7�h���L�=�w`E�^�b���md*r��l���\��ә�[�cm��ϴ;_���eR���B K�+������%�]��+Ҟ����(Ĥ����s� ϞIn���c�����1�
�acm���?n��o0b��<*�g�ض��'����XyV+e^��9�|G���x+,�nP�S9��+0��?��fߝ�Yy9�����^A��v���������,��_����X?5�� Otn���It�H`K��s��Z�Qd)�J�1l-�vy�d�
soi_d`(�մ���u32�<��_��n���'9Ēn���{L�&Y� � 6����4,)�4��۲6`LP P�%ߞ��ʦ���,��%���q��T���3���/1�3��g.�s���5N�9�Ű�?���v��L�H�6N�ϭ����@;􍋏��W���Ћ~�x(D=ո��.{d�z�tYL�rC���G&�j�,ug
�0��q�����
־�;��<#;�X�V�D[�[��[46o<94��Y4�f���l@�H;��p���nrd{�c���l		Ef�#Op�GVsD���.WE����.�t�������Q��S�-��|_It#RE�#�n��bI��6�|�Yv6r�&�O5�Rh�i3��c{=$o�t��r7��.�w������Y��D7��l���WZ��E�.��� u�{�]̿%��q5]�Џ1N��$+9�f��?|�Y�'7DN2�gK>kXX����2V�q��/:ܜv-h��Kg���H1<�>A��Õ�1R�O���˚`�Yk<ᝦ|��\z���LA��x?r"��T�7��y2s�У��T�h?��EW�[��/ghX��!�閌��5J"��A�!�$#]:�r�0R+�bٻEt-��p�59F�}�Ϗ��������cco>k��R<O(,�o���ˑ(�X����l��.��>r̻d�@��i[%����)f��s���m���^n��j1��u���B�9Z����5u}��^��@fG��'�_�:u(2<�_w����G|�р�Z���w�`�1�#��j��b���əZ��C��Ag��O& �����p<���D@7j�)Ж5�r>��wf�ʵ>%	�b�jz��y�>�7e�c�@V��!��y|Vw�$0?�b���-��=�mbp���+r&?&����D���ʿ�X_T�;�!݈͜�U^A[/�W�����,Y�k��=ٮҌ�IYwc�v(��a�\���+
hFTi�)�;a4�X����O�Q�����"��ET�2�%��d�a� ���֪����r=�N�_
�3�_>�F��Mq������wy�ҡ�'�dBIӆ\��U��
���?q���u�R�5i��x�"�V�H+�
p����/�5�G�x�[L8���W����混\ʖC*�3�(�*�C�ve2�������뻜��,�tJ�3kWG��m�"��!�K����Y��1���9qSU��L��-��Is�1�K��~��]��p�Q&a��gБ�~��w�����)���W�J@71�x;� �RK�{rXѣ/��."F"�V�����GZ6f}����qK�����o|�:��ϼ�X��-��WۂzpE�w(����Ɣ��V�I��J�v�cg�M�ݎ���_<�C ��N��|ϋW!�[+�_X�+�����$!P�Y��%Ӄ�m���@Qek9u�z8>�'=|�BVK�c`c��������T?S�b	�������J?���D��G�qBK�n��gm�v~�f�g	"OT���5��g���v����d�DWf�f��F��d��8�_��|�r��L�;�B⁝_�WB�{��R��9��3�����~���ׅ��ۍ��,�yϫ�֣8�e�Ѣ�|����]d�n���_J��Ed�/���2���(��7K��e�BQ�W�A+�K�(�b�n��G�Y��)����������6��|E��
m�����|BJ#�.Y�௜������:{2���u'����t����74|E�GBM��v�wS�,}��yS�����m���QF
*R-|�?�SكS��۫��AĬ�7�A��˝��$xٲp����X�0��6D��y&K;��T�p��:�r7h=)Tv�?^�%��3˷Ž
JK�	���E�;u4wK\��d|�B���|���$9�-��{��ذ�g����Wc�#�ԇ���\;��y6?	����h���>�c���#�OJ�C��|9��;_IV�l�m��ܟ��S<p�c�ںz���G�5��p��A+���Zp:��o/ߙ���e�H�Դԙ�����n)"�i咯J��D����)��~~�W����8��.Q����0�Eo�׏=et�κ���q,$+�)v����ce�J9��/5����V.�0����wqR��%}�[NHɲM�_˾/&�ޢ�L<�z���G&
��Sg~9���P��X�H�K����M�R�GЕ�{�[|,^�obi@J���]{��t.�h|;2��~�F�9tnsIRuk�w5�	"���c���K�Ƚ*��{�}���uRM��CcxB~&}mJ{֔��'pS�z�b���l�O�Xa�Z��vp�纻l��m;���K�R�֠�h�_Ϝ+1���W������-~G'V}��Y��b�~/1���,�Gv�f��5��$�{�ə^�s��5�µ�b��G��+��A����D�R�W����=���������ݵ=�;S�/K��DpmM���7^�:���{~J��9 ���O�4�*����W�\փ7����SӹR�Ɂ&XcP@���UW6�� q-z�#��=?0���[Ra&?s��3Ȋ�4�����X�G�$���>�"�;Z�����8�\�h,WGWؔ�$}��mΑиy� �P�5n��]#;�I�L٫��=Zym/yc���h�ъ����_��A��W��Yu��/�uÔB�ʷHgX}�kE����,��v�fk,m����UʡnB���֭�}�=b\g2���!Js+H�vL;¤O��ZK�-��_#��g�?�DڏPS��D��<�>f���g��K��K����%�&�܎������2cj[��F���mأ[ }̢�DE8�>��/��2����K�o��;5ȅ��-/���֞\Gx��P)i��;�;��Bm��#Oz��<_&�^:c��#$�N�KZ��T�u%�n��^7��4�[Ib/�0J�?lg���YY�?��un%Z�"zN�y�*���gBFGy �x�8���y(�c�ԭ{]������$Ez���,-��2uO����Ԗ����z������ͭ�2�|f.�!�0��C�-�ŭ�OՖy7���Y�m	�47���s��~KL7J�xJmw|\��N=�������(��}��P� σ7;�^43*�j�Z�EHфzDXj�����h�\� ����hH`d�"�L�}'GIS1�
��~��+U'<�vz���K��h��?Sp��O;ig�B�&{�e�z"%5����b,T�!eny�B��n'�F�x�*�Dq�����Y�E� f�6�õ9>7c��8�
�7�IODUu�����x�^,�I�N�T����Sa0��E̛&��˩!�0�'T"��/��|�����2m�?SJ�z��XL̵4b�޶ݡ0�Z?�m�;!c|��eW����&۸*�t�|oo���c� w}�~�8����<��b�Ei�C܄IO�Dߔ�_w3����<�}�~� �L��3�qY+���TP]*?a��~�>S�냳)�A;��$�^H�v��>/�ft�bU �-��iWٽu��* ~GjRs�X����Ğ`�Ocv&�F|�N픵��ut_Hq���7���7MFoG��#���7�=��)F�}r�s�3+������Q����qU՗(���V��Π�DS�V��
��w�ė2(KQ��BY�6�e@�z�h`ۖ�����q(}����� �r�އGQ9"�
�������0� "�C"�C�
JJ��P�=��HK�Н�~P����?��\Gq�yv�u��ޱ���@w�O�0��!e�դ�x)�� �%����~G�m+SֿcD�)ǒVZvԔ�*t����Ė��h��%�z�\�gp�α�������L?©�5}~��~����Ǟ�f�)�L03aݗ-�n�':��"�"$����n���U��:y�5\��a<ܳ&�y=���t�c�ܮ��KJ)B�
l}����ģ��k�D{{s�h�?>��ͧN�h����/e�0�t�Wa�󔨟���,�,LU��`���"5�Wq��m5��v�]���Kh���r%U3�Т��6ZQ���x5�Ek��Q�<3S�e�\�A<���n*3�	�t	�t${N^)Z����K9[髠[|���SeN��+�N9�&��f�Cts������O��;r���z��pFL'55GY_y|���������2%e��ק$��33Un<]n�	{"%�$�x䢭�x�sr����²(q䬯���F�ECfD�wh�W��F��e+��馧���mp4�~X���2(��;��n��'���?���y黓�{�����9*ˏ���D�DD�?��~=y���ۮ�R7N�|�#���_[g�˧�t�>�m$'�h�u�*G�F��tZ�!*a}�.����N��sŀgޣ��s_%}|�t�Xӿ�ݩ��Ԓ}���(��b�#���k�b-lY���j]���{-��iO�$���'6���-��������ȕ7k�9��ST�6o�#^}�67�֪��	�QU�JZKE�N^̃�X��앖י$a>P`ZXT�=��E�!$*
��"��u[okk{�
�����O��|�Z﹞t��d_�9���������ʗ�d�	d�� O�RSM���<Gax��X��l���� ������)6�?!�����h�η3;�͆�<�g��8V��qV�*��n���R�^����OO�~�N�G���4識�	�����]p@C�4��>W�`���;g;'>�ꙑ�J�!RIv�rJ_�5߇,^��-�KEdk�ol��Ő�_na7��2?�w��"��gG1%%%��8�F���S+���ȣ��67��糐,Yʆ偗����#��E۪�;�g�T�
���4t]�jڵU'�Q^�T:y�Ŏ<�nw�ל��k1��%�1GA�=s��r|}O?n��C�����������E:H��RƊ9�EO|=龿�;^�:�o3����xW�,�\wg����t*��cU�!����r�;ꍯM1L�йp�d�X��ϞV��v}p�������$��3.r�,&�h�숖�ꋲ-��7��z_m2�1�p�e]#�y��Žm��P���[�����ѿ����H�n�@���[����U̐٬��2����M����~��]g��L��z�;��c�xZ�|��Bx���{����m�$F8'��"�a/���no���ew���C�����@��aə�H�=�����{O�vT:�dcg�K�i�$��z��qKJu��Q���)�@b�С�T��B�p�h%v��:e^o�zΛ�J��ի�g������99�����i5�����g3126�x���{8_p��8�:LG�^:�ly��ezBpo����z��Tf�2_� �}�rm�D~̩nS.��㣍�X�C��P�1��-Z�n�g��v�x��:.�|�bΔS��fOr/���SU�q�	�癤�Aq��2��j;�w֣���6:kI�3��1�8����ڶ0(bQ��4?_�j������B�?�GG7�bg����pw�t^"nV�1Gm�v6����i��W-p�:����UG��l�߫x/XK%����|�;}��Ā��iB��FP
I%�J�j��K����o��HZ���9�N��s�MJ�oX�'��^N%��52����ٟ>]y��5��ٳg�deU���P�J��e*1�󽳝I� �����}%�膙z��N3nͩ�vF1k�YE1��dnH�e���R��T�z��~�؁�����VlG��D����:���X��[�x���tFW�L�s�q�b��MwC���܂$��c=����W��������xQMc=_mix�:+.-6�m�߽���|_�f�-�Vz)))��ϒ.s�ƨN�(?�f��$����l��G�s.���p*dp������߿:r)|���Q�]"(4WUQ!ϭ<�0"S��.de9�O��up��V�$i~�H��xW�QL�~7BG�Y/���Տ����j?z�X+F~�����+��\c�'A9�A-�����5��pB�^�3[��p!\��R0$�|VVpe��
���)*OM_i�2W����8�&$̬˲xn��z�j���q-&뤊㐰�.v��k݈����{̓���;�B���;�~f�U���.]�R������⒒k�q.�S	���XM��@C�]dӆSf�ˉ���Z	OxE2�ߗQԽ:���x6��5\z[h'�j4_b{�.
�O��ʦBBXs�:+��>g��V�Z�ІN���H����zO��E  �
W�"̨!�I[�g�;}��1���������&(6�����t����Ԫֱ6�����i�Si��L|��U�9�
�z�06x�����!�e-�������#�l7͠��5`'�\���5�{Xoc��;N���W�i�SSщ�5�#I�p�_�Dn]��''�=/}Æ'���Q���M�X����r��D M�q)��,���������$���h��̿��+)(���w;��I�5G>IUԷ�*hI�_�G�j�:��MR:NTy |���f{�q���M��WMM��[_����<�<łh��ݪ4Bn��e�u>����	.]xC##3vv����H];�#+���`AAI���@GG�x��C������V��s*UP�II���Ϧ�)�S��[��54"���B����з�" �@׬e#�z\���Cm�*��߼�E�
@�"����"5es�g�!�zg�ݴI��Qzy�L�rv��͛*e`�NN�5��t&5X�k��̏�/��(��#�a�T:�a��2F#��V'����}������ԉ~� �ڝV��\a�S�� ��7��4���֚�(}��e�g~�JKKsVB���F*J�5\\\
����r��[B�{i�h�GN{ss���`�^�����(��껲�&�q���Ї''0ؙ�i(������Z�,���	n���8�,�|�ljr�\J����6�(����lj'�<|v������8���g�1ek����w��^h;��?>�EşS��aa��H]'H����g�J
��mJ�|�F)x��\�\s�=�T��"��>&�yn��s�����^=*�?�IFKkonkˮ�#�l-�|	�ϢUt*S�ߴ�N��zff���`�i��Y�MLL�i�E�Z����1}oK8�>_�3�:��g-�o2���µ�YK��,@�m���U'��C!���Ly�X�)H*.�P:�^���X͛�����C��tez�� ���.S���F�Ħ7)-�Om`�,�iM�I�c��d�l/e�T��G���$֟�n��7o
a�ast��IϞ�e솲_Co�p��qy@�ϫ���� Mpʔ�٥[���Yw�@̇t~P�����4E*~�����N�/{�+9�))��};�P�`0�DK'.0ޕ�.���q��)ڙ��Sf?�>Xמ�t�̃Q��l��Š�)@���m��5����U��Q��L��?B�.��r��Ȥ�.��\�%[sNŭ���=J&���
*z.pgCqqqӃ�U*n��v	t���s|�3�ɝ�d?�'�蘘�eW�I鸭�A�.
���`�fS�����D(��Jj�yp��6�?"]�e+���p=	�X�'�ɰ�)�٩|e<+y+�5��l ���m�U��[i\��V�DIu{���b�'��J��m�5���T����Л�q����έ�������>�G����6���8�h��"X���gɠ�]�Q<�>��٫���[=��{x]�P9֊Q�n�'�D�`sX��]�#��OS�2� &���	]	;i+q�L�N�Y�0�I�-8s{�f%�;�l-�gt=4d��:�����n#␕=��L�S�-_��݋�}��Ĕ;0�=��jA�MN}C�9U�#�th�(cy0�$,�}���eK`aӅdq ���d�B����_K��k;B�ef�+74)g=�S�H0W^�)����PϠs���,��W�AF�;f?{���2J@���r��{���g���od������ȶ����Bw�N��u��-��<���X6NH:�Ƣu����㊓*�cI,�I��F$+�_���L]�vH��˚w������R�G�JO��(�D;G' ���B�#t+L����ǏD$$��6_@�X;G���ܬ�CQ�y��F)���<���L��6g�1ܘ]-��&�_��`,�z�;V3\�Np]*� l|����I	 7M*2==�e.9���T�],����`�u=������D�=��w���:���R���u�Jlly�E>h?��&��o����y'�����X�Q^��7�v�^rY����xql�k���� ���QRA!�>�!�4�=�!(

��B�$+�סZR����e�*�k�
�������y[[����@�dC �2~�h_����	����e�&��P.l�h^ņ@���ii�j9���/Y�v��a�L@�2�����g-∁
	A��~�e������Nl>r{��)4bU<����Y���-͈&��a����#��]'�PS4�j�f�o�U�>��o��e�ͩ|5"!a��8���w��SOp�Ƃu߆BhF.��~��G���;Tj�������OxC��I~^^Hh�q��h>�V��ݦ��ϣ�Q�۷Š��s����G�gA(�L9���}��0e>�t� J�W<�TW���f���������@)�#��à��#�TPQ	i�����k���4���$��c�<��y�����H�e�QU;7����{����4h&��8�o���������z$0��F���~,�3�|>Z�?�c�w��Mff�s��uҺ�(\\�|0�$���X�X4]
������'�.�N뾡hYw�ﰥ����wƵBJv�����%^{i��O�����D���;�?~�o�v�A�J�a���m[�0�����n�.w��>�<��./����Yٗ�5�ώ��*֒��	U�xEH�t<�oM�[E����eF̹��
�M:m�$�nR3g��������9ם�O2�v�@��I�y���l�_��'#�A��&��A9j>E˺��K#�aoߺ7C5ej�;��?��V�4:������o�Q��"z�||@�� �`&��:�����	a�}��B<p�^������N��ged�EEEe����8w&<�O7��f;b���� %]Lc���puv�m�uo�(P�#�디�������c��^t��ӭ\Og:ߗ�WP8<UhgkUs�\�9�(D����/pT�����歳���Z��rX�����Ǩ�E~�����Jy���n�e�6�9���,x>V�$������/ĭ.��(_��X��%��p�[m�.�U�����c���ɐ^EFj�H�9�,�������//���:��(�0i%%%R჎���V%/l])�]�»ahr�f��f�z���A����2s �333+��������4⺜�(� � %������0l����C��T�n�Ny���0=��(�vg.���j/n����z�g�O�r��JHH�W�k�҅��bE+BG^
�ꯡn)R�6�O`���J*�:	�l�C)� ���>�~Ip�x�oݥ��f*�����N_�#������UH����d+]69b�7{�;�\����i�����B��j� ��I��K]3-��_���a�m="н��XHt����٫�9(��y�c"��r����P�'vQ���O�7�g~c��:W� ���Q��&�<�lh���3��@�#cG������O]�<,ii+|�������ի�1.w\�n�"(��ǹ%��ޝ
�]�^=�� ��͆�H8;;;�� P3��E�����Rn�̠5�;&���'�_�*:�}���~��Ya𘘒2�>F�?zA�x������(Y7\��}A kX��Y$4����3va��P��3�����D?ck�>_������, �O���������l&���lb�����6�	��?���'$$t�z��7��B�I�7����?g�`�v��ω���'���+�ڿL�O��w<z��UlUu�����&�ݻ ��!uEP��!�����"���KG��	@AG��v���!��v`�@W�����K ��=555��V��z}7��p�&�����ng���;�2�IL�խ��6٩�t�?�"6��>�e�)�\���kޯ�W��'����^I��~��Z%m�L,�5K3������W���x���Gh`7 �e �)��莾2#Ϊcp���fLh(�	+����d�p����֜��H%�N�y1@i��OC���\����{(d?����o߾�Jw\�p���`bb�����+J�?~�C�5E&^��]P��0�Gy-NDU:�g���ݲ�
����U�T$%�]fվ�������2�R���D��ds��e���A��o?�@��C������Sh��Flq�;���Y*��ۂ���VW� �I����4cFc�{��A��ցG��_�N4L�:��àZ�ȏ���Y�'r�h����\s4�V��?O���J�ҧ���> B*��c�A{O��H�Ha�*��T� +A��ai��(҇q2�͛�j"���|�N�2v��Ȩo�
4N��v�0��}�t��v���<M��o��u�_��G�c܎0�-�2C�Wy�gf����C?e��)gBȞ���峀ׅ&���E�9n@s�|]|λ�A��Y+��޽���-Y��+�������R�Ӝ�Ν��
�Ќ��؁��1{xV��!Tn/>�w��ֆ�
x���E��ԗM�m*�?�0n[
�2ƕ����H�D��Ѥd�9���c�h�Z/Vd+kQK]���L.��5�P��}�9pô�.�I��N��{�bon/��K���R�(fm����en5��!M���Y��$���PE�]�!�}�����:g2�455��@:�A��~�>H}Wl��T���ru�������B�	�`��:V��G|jS��c�@s=0�mk�q��2����Vk-bz}�0�o��$pQ�æe�+d.0/��w�Jcݓ$�嵜;!�ԙ]v��PQ��,�p�A�"��%iY��ǼO���:ϫ���?�o���?�N�Z����AiD:�cR�?}��9�������	�)d<6�4b6	��`��);۱A�>�^�ΔT_o�/PE����Ў�,%�g��N;�_�-<���k�(=g��4�Y�*Ğ?��͛N�ԄQ��{��/�J�&���ګ�?�F��-Gӿ�W�ɮ�ʟ�t�`m@����F�������2�33�����-��Ш(s8t��Kr�0�袬Ũ�H38��FZ; �Ƞ �	#�"S`8�w{�Z��s_$���`�J��)����G�Y������^a��S���RJJj����-'�δ��I�����3��MEG_��(wX̨���u�ɝ�1��(S����|�fN
�����MvҊ	�گ���58�i�<l���>�����i�9��/ t���c��|�r�s��K�!��d|jk�_� �g9��.����:;`N�TGc>�2��aa�	�ouuP`J��e�L��O�s������ϼ�g�8�v���.Jq��w�u���#��I����󞧷����Yj7C%�&y�I@�XRRו,��o�,UE�7�����޽{?]U���S�y�ڀv�_�D���c}���YYFF)�l�������y��h�k�N+�k��U��,���Z��Q����J�����+˥'a^����#%�v�Z0��B�.��B��1��3� (��ǁlLL]�g�i9�d@�����:��2��׀���X�q���M�$s�7���nb��T�%e�Mt`�d�9|0���8��<�hg��o6U��3wbJ_#B ~�Lo��a�1L�Z��B�_�f�&�G�4VH������[��������x�v�ܷ4b���9c �̫�o���՜c�\�ǹ���� UJV6k�z*ݝ;P}� �k�Sd{�$H)()��h<S'��0�m��N^T1��2M�}���cL�n�U̜��'I0 �CK�s�y�$�
~���t[V�}��"q�g`��(�щ�V��������%�t�C���B^���{#|w�e���p�M\/*l����)���£�1Vesw���`MH$5Km�M���y�.!�͞�7�0h	��ߺ����W�L�r���s�n�J������˓q�++�ec��R�vXǈ�?_��V*Э/��h���k������j2��=�Q�툶���B�O������m��^��k-y|1,�-E�QӼ��n�"�ksp�l%v�5q�Ń?[�T			PY[T3K�N�R������M2���-��>����l�K]	�UK�@e�(+>^dnn.e��Y�gI��^'0�J<ʬ�3�oM-2 0g���}������m;��)k�h���i�[�k�������kx�Mb��с�����d#�^3�6ו5T��=��H��5
�b5��+�{��;}�˯��֋���S�(����1Y?��UTټ�R�I�D�YX��0<q�q�\�n�|eS�Y��M?��^��0=<�E�,H4�bI��Yu�v���YF��(��r��o�/�(�Y:�=.�+d\�(Զ��.��X��C��^��Ք�>�9h�2ٮk���ߖa[�W�U�+��Qop��U�VT-s�2e��B�r�՜�=���&������n�O�Q{l��r��c+W��e�D.���z#�Z e�܈<D�
��J��2�A˾����-dgX�Un�:�3.��ܮ�t��!X�&�$>��<2b>��'`���ޘ�^r��$��+	Ə���ѣ���i4�,x�8%�))�1���n���P��G�?r�^�V�A_�iǂ���;�5�%lv����R���i��A�L���vV����xI��{��ݻ����-�5o|% e�Us�E'��>h�3�<���k�������w���|vnm�<QPN�B@Z�0y�?�
������5_��G/�t�@�DBe���0�{�q��M��xh1���9U$����6Oq]*mXUlH��i�}�a&;�@��#&o�8ם:o��w<��я߬��U�y�6UZ���=t��+����g�l[����I�2��u��3��}M��T��*�g�[�*�RD��i��V%cg�R-��/��z�QY���wA��}���Ơeh���5>%�E1��3m1R��h�> X��q�EP*d�V �!�n(�;�[���˗��8&;��^t��;�NP�)�� @4����񵚝�~��2
@���DF
��[��aa�tڛ�����T�<e?���\�)�ں"�&~��T�faׇ�bP�%&!��e;���B�;��A�YP�N`?B3��C��M��9T�����9X��
���hTSQ	�8PI���;О1�������m���@�4дR22*��/�z� �7��>�:�B�6���3qK��wZ�\��R,U��ٗkjB;�*����ʵ��j���
L�d�,xL/�SYo�o���E���^$���M��RoL��!o�R�6"̫_�>Ѹ����R���9��wo�v�0r�����(D"ev֤ФST��~���6t�locζ4Áy<Z*�b��J����Y��hO�he�A�29�22=��
�B#��CJ{8�\�l��p��T9}f�p�ט�Sx��;72�>��i�|��l`��鿦�����%��aHT:o(���Bu��kNe�cY19�22-9��{1�>�p�'t�ǘѪ7?/4:~�Lù���jO�Y�u� >��4A�p^���;:H�U,0鼥�4�*`���t)�P5�a�(s�b��YfT��P��٤�=績LN��25]G*�G�S�b2F؎�0*����_,���v�r|�����L��] ;,�D�<��/�y��k�9�
��q��/�9�\��=	b� ���K�Y�E��04Bn�kx���?F���O(,]p=��ۇ��.N�6
�*.2Q9��ʑ��T �A�.�p������=���U�g�� �P���k���C �鹹�O�c��	Pt�v^���NVU݁��f_c0=�����!L�)ɦ �4��	iU �&"�;��J@q&Lmu������R;�[K��(���S���`d��
 �z������a|��}��M�Ѝr9dԮ�E7&�r�#oc�bX���fYW�>�RE��x{cg"p.D�^DM��qM��E _�XF��["8Q��=&1MN����� @����o�/��A��=\��@� ;�K5�o�L��E_rTL*�#�o��T�*�q�[�`0�P:h�\��`�*�1;��j�Wm�����U(6@e�U�0��ZOmfDf��fgg������#�z/��c�V�].��	�҄	��h��lS]؄�b,�����9y�*����3�/%Ezf�h& 4�|���+�<�v��_K��� .'��v(�2�"2���eR@Ũ Ce��14�͢[���;]9գ0;'xho������:��������x(�4fUn���j����-Sggg(9T:Iի
�QeLmm-5��\p�����d�� M{���	b>��]�9��<Pu �T��ǥ�c��@Ȟ��A l��$��1Pq�M`|�I�����L�R�����к���F�U��Gt
*��:��Uĭ=�hk[J)+:�W���Ⴌ��v���#��f:���a�m��ƒ��.W��~�h8��j��%��y�J��[�P�\(k�p���]����K�h}�fC��2&e��QK��m
��A>Z��k^�`�M����C�'��Z�^�>BM[ۼ2����4�4q��О҂CyMM�������[�/3ݾ-Dx��'�a<P>r(��?~\s�P	(��B�CCCT˝�v���κi�$��F1ݙl�?��秪����"ch``$^�ZB`��
j��� #77`�Νn�4����~�?_��v����̵��� �==N�>��ֆ���&~Qߠ��`����+n�����"�W�� ���r��5*�eZkL�C��!�â0y��.�d|���h��R��Y�_������� �Q�V��J�qE�������Y�*��"��s�C'���~��U�H�C��*�W� n]eu�ǥ���hXI/(P� �}|n��dK_�r���u�sۋ�8��]�z��NE`#ж��L��j��������2���<=!65|��y��wd��PH�8<Tx	�څ�{���'x�6����}��!�×P^�tT�w��M��Ha�%+�פT?��搛i��6��7��_�1`0�j��x�����6_jλ�>?�#��k�(�/3��]��{���FO�Ӫ>Y��<��vc}G6l�G��0�J-#s���X��w��?�}�\C��iK��\L�Er���i�%e�>ǐ�2ұo0��_�S�̞t`��gA�J��H%n�E�TЁS�N4T�*��a�@�k Q�o��N��11��Y��񖆖�k�����AfS��iN󤜙!�xU��_�a^fІBf{(�x���F��5�����X�ɦ���x�u�E�69�&�KF�[���y�9]JS�u���1~r��1Ẇ,�v�I_n�jg�O?2~-��;�5���}����U�>i
�6�պb���D�;�z�UA�˹�sf��I���?&Z,�6����y�b�3?��[�~ H>yu�;�MI����y�(�}��Q�k����)�NI@���4�,��г�������<��s�I��p�x��ICp���>��������A��ar��c��C"�0FgA�ѕ�D=�*�/��H��>R-XL^;?���8�[q�'��R��~N��~$j��9�_6o��<�"���a+5V.���-?IB��_Ŵ��"z�=������t<��Ϙ����N]��(��V ok�/ū�"B�&����Z?�m��g�jJ ?��ǽ'@q�<��Hc�3��m+���y��fL�C[��rx�T�yʚ%z#Sz��3����1�^fp�o�=p(\xӐ@��G�Y�$n�!��`��9CF�u���~]* $mHtt�y�5���e���h1�f�\��l�8�v��ȹ����S��Y�p�}��KT��I��qDk��D�m4?bjا�<_��������ע�Q_G4Z��Q���s�[I��S|m嚆�>��w���Nk�J�[kf�]��D��PѸV߯��IL��P��D���QjҜ��z.�Vh��UuY�'��TB�hR;�ghC��E�젇dǻO W�Oga�z��F��lV(��c4DZnqM�:��oXD�~�ǒ��+��Ъ����y��*�W���GU��mu!Ӣ��]1�/���|�f��b���w�Y:qx7�+�NR����{
���LU�QZPO���f7���^	�y<[+O�b����zy7�z�|1�U6�bE'�G֜_V�/>r�����m��y�y���qc����L7�� ���j1T?���]�{�ȯޢ�1J�1W�� v�a^u2�^�Z�%}��k̖i:_��}ON<|���B�Z������8��z���c�:GQ�]�e�Nt���O:�
�Zk5�T���_�{�u����[��\�IةG?�b�4�	��δ082X��Թq�zn� �t�����^�ӂ]ب����=<��꣮��sng�|�(�D�'�Tb� QT�ۿ����\E}�U��S���,�� ������3=L$XP�<����'_����RĨ�t�Ǯ��*>��T���|]�[@��Bh���c_A>D}��]	�ˡ;�:D|a�(r��������|�G�A�h ������\*Z6�ˊfLJ�1�I$Uл�����+#]Ӡ��EK���'j$Ga0�7�Ȝ���+ оta8��l�fP��%�$�˃�ٳ�����zk��?gV��Q�zN��R�|x{�GS�)]J����@����[QI_���z�?���e�H�>7���!��k��(0�Bz�'��?-���/?,>[ܣP�>5�~楿��J }��-!,~�oϓ���NI�r��O}Y���aS���Yk�?m���O]0���g�����Z�&>`\�e4��C����W��~��<�w@���T��z�$y�G�⨵p�̀gj<��ǻ�B�l�Wg��5��&b03��jk��i���#��	>VS�'� �go����&vb�m�Wy� �C������WF���ܯ�h���QN�7����2�%�l���hМ&Q�,R�b���z��v�OL�G�vJE{O9�2&ND��j�"r3����~>��H���^{7�j���^���Pw����:HBП ����������8�`t�vA���/�Gw�B80#\�B�^p�3;u�[�ߨ͠#0�~H���z�Y�B��*l��h���$��Z'vdr�9NA��#�z��\q�$����a�p-��u�G:$���F�)���[�,�0��h�ӄ����ux%�+���w�k�A�OSXh`;�eq|��/���c#q�������W�g�d�S;���3��i8�.��n��jY�}b�)B�b��Ӿ�U����ζ�"��4�7�_�eIO+���E|
<d����לG�EO��5�#�����ݖ�^p�}e@��Qc�
>�;q������ω�tI����D��xi|�Wʀ`D�ԎA:���?F�fi�|d�}O�&4}�<u5�ͯ���� �S@m�R�Z������K�_~ =�(���4�J&x�1�Cs���"O�n޼s��HPr���1��p:��t��6/8k��b��/9~�l:�D���k؋;��7FPK�#��wB�T�p�3�nn����`��%�e�sLa'�8�Ϝ�`�+��b�r���4�A�If������[���,B������ݡh�է*£���ܦ��ϖӕ�����>;�u&=��ԙ����D%���M�v���o���G������_8҅��y&�}����-/���؇�O��MZ�F?�dk-;c
�_��.S{�|���=?�
5�Dǫ���u|v����v��(ce���p���0�/��a?JL�����J�6e,�<f��Ӛ�nT�O�x�{5�6~.-����o��d���B����4=(w7ۍb�-
�*E?�Y��|O0���V�+t���*1!��]�O
]�ʈދ�)��aޙ�V�]Jo��z�����75_���l��}�3�N�D"�Wv>_��0&�B�P6�g�����<90$�%�2D�R
�5!/p�H^
�3����|�S�����3����LMer�	�q�k�_�]Q~�2۩1�����k�9�g00��eb�g��l+ѧX��_�MBmt�AT�힏G�.�K����?V�n9>:3s���^cV.�禾8�w���>:zo��#�i�����0�3����_��H���U�t�9�����['>G�\���Ύ����K�{鳋x��.[�GnܦV��ic7�Q����3h�+oB�H��t |�m	>%j<�v�k�ve���x�[�������|ܲ�n}��-��5#U�~�K5C!��9�ش9����;�y�=z����L�u좍SAQ�--�EA�Q���0�J�?n�u��9��Ao`t4=�3%�q�8�%j�@�x$�*�g]i-ͭxZ��������pƩ����������"�݌���&5Ra�dN�[B����Fu�I�o��]R���VfX,̸z�Oji��oڭ�h�-r��|��"�s�����}�E����B��~4��3EcϽ�s_��\���{
ҚB�W�D����ϴ
�/
y2x�IΧG�K��j�3��Jta�Q�^M3�6�u���q�("��P�n�����-M5�%�6�˷�&?韙�ĽҞ�|�;��ׯ�5T����2�u�P��ݷ��Ԯ=�t[����X��V��_o�� _.ճI_w�^��Y=M�PU�e��������QHu�Px�>BQ-t0�"�����9rYZw�4��oThWI��ʼO�Bg~9O�77��n8暵~>_��L���nf}��SQ���^UXK�z��κ������{�dɦ�;Qj�	��m�F�C{U�~J�/m������IEtl���3����6�k�/7(�����Q-q�i���TZW+e��"Km|�]�΅�窅[�߭�c�x����=ףlvn�Ĝ��+=rc]�Lea���6F�g"'���/���
U�o�V���ی�g��z8�RN�v�`*�A.�,��j[L^�͔Xg_''L��xmv�i;Ayb�α��CѦ���q�[
&�żQ���8n�pt/��[��o���I�؁������w�����/���Q���1e�]=z��D��:�#������5��j���~\W<j#"���4!�_$�����[B?�{�c����'�y�V�<h�µ?Ͻ�����Ҽ�	���G�<�;r�q��7��������y/�<�>+�wm�R�-��F{<��u���$ò�e(���Vvu��� �v>�z��Οq��� �}빷�	$��DsR]�5�kb�y ���w��$w���,\]�d���ov�e;a7I%n�,�����2�Eƴ��x���	J.Ҏ 7�Rv&e�	��V�����G�S�ۺ�j�� !��,�xg�?�� �<1�����FFTM���褍�h���?|�����a��.�%�ݕ�F�M�\�R�c��h�����}1v��͌v%{��9n�E�!�͑���F1O�b=�_�E���˻݂^mb���߭psY-�%�pVAF�n�}վ?t���кGuv����9n�gr��e���<�Ke�M�g�(�<o�uվ�e�d1�FU�F�w�+���#k��#�cx�c�O�vo�ޯg����w �R�FD+~��/��{�	4�Kr��:�=��8�Y�s�gB��5�3��EO�Uj�},o^:c�{����N�$���k~&����xDA�'�Fn����M��S#�����Ky�#��V?N�+�B[Ԏ����"rt�`ZB׶�Ү<H4*�!���.�p�i��V.��l����T��g:48�~�2d�K��%o8�2���;qDe�ly��3������g�6�����JK�2w;7�D2P��Z��c����v��w�����D#���8�`=y@7�66�8��5$HN��!rA������]�`�`�%���73| �*n���@Ӭˤ��Ye��.7��?����h�1�����`�>�h��ے�Ͻ��K>K�<#�=N�C���O�a�J��[&f��(��,�ן*���2ɚp%I��1n�P{��6�U7;��R��.�}���d�?��7~�x�#P8�q�м`goY��~g��y�(��.���:�k�d�%���:X� �7�t�ZO&�)�'��/׽8r�8��t���6G�7�`���Xx�}NQ�,;X��!���lg���8�������٣����������S��4[��Qr��nK}��_3ދ��t�P���y���RΣ�#hr"8���]�������wul�>�4�f��.y�X��} ��{XRY��+�\�g�RY�Ԗ�a���Vr���	0<_W�]�ʒO��`ҩp��{�l��z�����llP��SR
���$�S?��W�w�����_��k�f���������Y��FܳepZ��AK�B}�5��t�YCN��%+�ym0�wq�m�*rnntWXXNrV�r�y���gI.nK)�U���d�,��
+m�z��=�GYH.	w��,X�S��$H3}�i݊�l���a
������Yƀ� {_�j�I���&��X�Y��x�����C��t�
)e�sc������խ��O�i<���	2���B��}��;7{�Q�6����v��څ��X��p�O��eGK�8R�<@��ѕXҙ�x�\�5���F��M}z�hƊ��-Yy�;=��TT<b���ե����j+��w\Qb� ̪� �=�7�w��6O}��G�]�3��}`a��$��`���,.tz������jֹ9߃zʼ6�ny��-���(ZSÅ��|��t��Ҧ#]����u{��l��5R#��7�3�7_���֭G<������Q9�n�-�V�b��)6�(҆��E|�|�^����붠rO���D櫻��7T*di:��M����,�����ſ��z�
(�x�AcK櫢�	��屟n~S>�j�7����cO�s㴶 ����Hi���v4O�;����[Y��`�f�-���6v��mvqjЇ�]��N�P�
� Ɵъҡ.�ع�d�dS8�'�g�#n��ir���h"�c�Y訲z�O�崁�ŀ���x�B]�������8\Y�"�:n[aa�mr�·���2~M��z(��ad�-���Ɠ��K��>2���������@Muk�Q���"M@DD���H��.�D���+��ދT� �t��Ѓ 5t����+��L�q���Ե����Dq���w�����f�͗���ML�L���� �b6_�}r)��ܼ�$i���Z�`{�&�>�2���V6��a*1mX�������-��V����}}9Rk�c ���~�M&���>@D`^�����S% _�����۾D�@g˿���6��`��o�^nn��m�<,Z��֧�fl�Qyfl���_+ALfj�6AɾP��-@� %�Vv�r�jv�]�0����Oh;~2�w�K�������uT�Y��6��}��qz�3X"
̼�_��+������<��k)�.׍�[߉��31�49[x-�����z@��%Ǜ3O,����>���c����n̾�)�e9R����l���1�"��u��ý ����,}����8������~��~dyv�ϢH���0�i@z/.0\��`/�t��WK�/�ڃFSd]� ��=?/��j��)'�J"������|4�1G N�1�8sȎd�������0����֤Sf[������,�bF>P�Q�m�t���E�_���1M��"@N权7�S��SR��Wm�ͭ����¯E�*����6;!a�w �����RF�Vğ]Za�
�&Eb]�Xaez��P��h����b�f���Y�����\y!���RU����R���D��n��d�OI�4��ծ�5ԍL���O7��8��nVy�=TI.�������O������)$����>	bylK�`}b�ȶ1k�#Y����	�>�Gg�n)���
���[?B�d��9������DgZ���D��?X(3�j����8��D��r���ݯ���LrpxU����!q��	b7�?��]jϠ]��V����E��G�~����˲D��JA��O����8��4GJx�_��V1F���[f��A���k[F� 	�G_4�S�--�.���+O����ٴ�S~g�%�Cς����@�����Y�����M�1�%F3���M<��W+DP%Z�����m���G"
&Dg��E��"���<��/˄sI�w�<�Iv!�?8���Oc�r5p$P9�겙�u(Тq�P��\N_���cd_p��:��:ъ�ݳ��;�r����8�s�Z�����R0�۝(W�������%k#������x�Ji}������Yb�x�+����3门5���o�j5���{�F�ub���A��V(����g���T��yfq����tt��^�A��#l����~�����z���Ϭ9	�n��
�"t���Qx�{ߣ����l��m��H=�w�#9z�����C�wD�)�|����ʼ�;��_�����1���Y��I�m�9$��|뾓׮olp����f��X �@r6�nI>w��¥*9o2�|����SN���jE���n�c-t�gX� ��F�l�1�o�i��6�u��6�m*�.��� ��"���ٹm������g���෈�<�k�ȝ7��P���Nz^�2�0(Ϙ�z�/�����ḅ�#pbӺ����/Ï�h$��>Nu�O��*���d��K�$�uüp��S�3;gm�-5S%��{;��G��䊱q�,%ƺQ,l�^��ϙ��\�f�~����e�q&����j{������zM](*�!AD��k�@e]����]�Ѿ�׶��?�ߘp�9#[�C�]��.-iSd��}�T�s���9���o�fFeD��Z�V	������oǕQڙ=����q�o�����<�	1ŐI�d/�VP��jS�Wո�r�F%l��z��/�%,�w�c�Ր�N��ON�pO���>���t5I�ɵ� 6�W�J`��6��]I���3�5�����-�צ�XA����2���?H§�����?r�]���j�@皘/��F��9]�]/�)c��'E�e޳,�\��`! ��J��x���ڸO���N_]��W=�8�S�.
�BT�\����<�������W�d�^~녺ףGWՔ1�w!n��$�aP��'yT���;$l��)g+mF����;sy�Dl���r�o*���uA�;ux��(�w���A�����"@a���	0ϭ������ ��e������g4�L� sTR�A|�	P�V�J[bzL����{�5+LzF�~�]�!�<N�I4T�'��l_v��	�;w�����%J}͌O�tܦ��w �� ?��+9gEe�@�A#wq���3�%
 zG�0C:���L�ē�|��+'Zl�KEتMV'��B����1Q�?P̯=�^�R<��V�>	��	��\��ܿ��8���"�vy���� ��Xw�#FT�J�?Ȅk߁55�J���r6h��Ђ��<��_�L_M��Q7Q���]�4��I]����6G
��!�%�N�0�ĩ�|��.����3��E�e
�`�R��31?��P0� �mAP�t��	+oA���I�mQJ&�����^uf�Y<����C�.. ,GW,Ӷ���-a���?��n�Q��]�buS��c��\�N]���1��0-����}�-gD]��4^��=�BV�uR�C��u��'؜\��z��YC�F~�K
0�d���X�6�67-��D9v�`8�<�k�KF�Z�{�7H1��k��ű�#�Ό=.�.!�$L�����'�:����ME�Q����ɲ�낕"���/��FD���.�(�1�V/1PFU�ץ��z��'�2(�`��MY㎝WG�OO�ț�1%��V�*�
��;V������fA�TP�$ى6ޙf ��`5ۄ��(��k�җ�9:� �/M���:=?J���ʵ!���B.�S��b/��f8� S؏Dw�pIW���?���7�sf"ց�`��`�\~����?c�ھ�Z�� ��P�r[Ɠ0G��M/�|��.�LY����=r��~���B�jN��*��A1RDN���*!h��&�`U�w�Km��& �&����1�D�+�V��/�X��NLg�r��֮�����Փ�͘���.
#����w`(� !�#��h)!�u>��&%�CZ'�<�Zk �Kr���It���C��h���N����eމl�&¡7�)V�n2�\D x7�41�`� �
MӀ����T��q�m��Aݐ��g`P��l�˺���}u�������U��'je�/L�]�p#I��͛el�=��hB4eY��[Vji��7�(S�%Ǻ�y!��U��,&�ƚ��|��@����[�������	���E�G��!Y�唇@��|T�>@k�L�z}3����aT�F���$��!�DP3���<q�^���.�oߕ�١��%w2�����z]*��3^��jw͞��2����=��N���h}X� ^�T�_��Yk�<��V~�bt=B����G����.a�Q���a�nģ��IH�.K��w�Y���s����E;�MEO�x���M��e[�R�>wc7��� g��&�����$8&*h,��ZoՎn".���m>�v�����Ug0��VK�nd�A��B��onv����-��sL�y�����η�
$C���C)F��W6�֕^����㱪�x�`�@F�m1���c��V6Ѭ�6||�}ϱ�K[Q�Ǿ�7����G�A{'��ktCf��{��� %���גվ��6�/H«P�3�����f�������79�@D��A̯*�_����ei`~c+���9���}�_2��u���˯~�IdÀj��טq���Z7����r=�[O���@Vht�u����&�8,���ϻ����C�m��Q_����0�3e��ru���+�~��P	y���E�i����l?�.�+e��g�Pa��v��j����2�Z�>`ҽa�hFJ�U�=��vР��K`�1I�48���8��v[ru�хL]�>�/��I�c9Z�`>r�j� �re������!��~��Є�09@��uC�a h��r�3�MgC�P0rE�r�H3t�ָEVT�vP���;fB�������Y����{|��z�u溪MHK費q�d�p.i������ʥ`��q1?b�*<��Z��o�����z��M��A�2uaJ�O�;�==�*�'��Ӭ��5��aKKߥ�ї����S�c�5.�����Փ��a��F���Ȭ΀R�����<ն��
�1BXHCH!
�9_�s ���sJJ}�O���JD��]���h2�9<s�J x����#2*�YD�2r�W塡t�VS�bba��DN�tsJ���ص���R�Ŀ���C�2�r�P`�I����AeE3��`�M��S��ԧ*�����z�D ��MJ�|�E<I"�i0A++r�I>nb�W`��;tA�L��u|���]��͡�⤝aȟv>�Ēg���S~��v�&�'���}r�n鏌�R����-��\�xRmh�����)��_����56G�L�-�7vح��C:���Lr`��K�J��5����OV��v���C�δ�f�3ej�������}b��3A����`ѩwŐ���R���T�S�6��MzԪ��Bb�va���%_�h����8B����ʤ�%v��)jhZ�������bb�zU<����P��0�]֎i��ee��+�y�c�un(ĸop�6�����:|�fw�'M�@}Vhܡ�Ս��a5�vW����M�%�{�=�%�������k��c�����|�W�p�����<U�����!ccf@�=i�Ӓ-!�;�?)z���[��V�?�G^����3���^�e�U��ۀ�B�0���U4j��j��^�0�5E�_�z���G�{����Ժ#K�tj� ���֑�.��c*qP���9��È���=+�:9�D �ȴ9_�ȴ�j(�����nMvhY�FN�V�6�/��sy��~3O_-�_�ڛqΘ]Z
AL�pwv��s���+�`�C �r��G�^��׍	�l��('կ�\6s��F�vj'��,�4�jT0��$\���b'�묖ҷ��?���m@/z}I�Fi4E�,G��V�.0$��C����ϛ0u�����6r�n�6Os��/U��"~x�ă��������Vp���MI���,\��Y&��:�&��C=�K����^ӧ�����@��+�4q�&����t����\ \��+Z�У�w��*�.��g����>�5m�N��k!b�o��:aM��lc��$@*����y��C��3��$���㜍���Vٞ��m���W�z�p���K�LV��s�{��'�&V�=� 6J���Jh��g(��/Y�"���	���N.��%Ѹ�
���m�`J��-\�<�`t�i���m�'�����'/�Yg���MȾʆ�פ�l�����Ax����b�X$|ʩ����d~0�Q��H]��j�i� af�"��ѹ�n�h���ݬ�M�A�w�&�C6.�4].ГX�5�ĥ�z�$�S�)��6�0�+A��O�Ϊz�c�j¥�Ϧ)�z�3���
�4�`t�r��7���SH��0����zD��V�2�����=��˥���]�R`ͱ�O���[�%�-5�E�{}%�Rð0����V`uB�z_nO��\��۷�Ć��>�"7[��;ۯ�K�{@\s���}w��7��w�y�k��O��/+b�s�W6���':����cx'z�)>�}�jpֳ-�%�Y^�`0�Q��<�@ �iZF��'sD��O�������L�B{���\��Ç�ԓ���~��7��SS����*���CK�w�]1�X�s��͕��L���Cױ�.\��LP���Þ���Ui���R�����M��ğS�ֵN�g�oکK��̘��ж��AڊW�{\����K��B���b��


�^U��?��wWޑN,�.�[`>.EY�Ӌ�$���'��C�S6M ���ͧ���#�@_�D���wS�$'m
[�F?q@W�39�Zr�뛝��o_��U��WL��V��^-O3���,-��ګﶗY^>Ї��;���,�u��%ꍤp�����z��yz�'�8�h����â��_k��ը$!�s�O���S7ט��966��f{�����/�x-�wq'������(nܣ#Z���M�E�5�GВ)QS����ᮙ�����h/y0p�Q�IȺz�t��b'���r_���Z��_X��3���}]�QÿӴF��c�;��ޱ'.�#�tu��P����̰�ML|,�b�c��5����p�{i�x����rH)R w�mz���q(�	�ső��������P������-�:=qZ=�[���T�>5�8�-�)y_�BA����8��`#���7�(<�x�V��4�|V7��؝<Y���M	D����Rt�ZZ���n��4xȠ�	���b�H��_f�E��k��L��.s�3�tl���?.�u���a�z�|H���$ 6m`/������u43_5t=
݋���4���O�r��&���`��s1ȰDጧ���~� ^�h�3�u����mΤ�g��y�4R��K�154-�уc���y�n�p���J��Ŏ� b(�{��l������9�#�}9���L��Zf#����D#R���`����p��r�Zf6~uh��7�/���&E���`��.@hy��}/��K��竂����ٴ��.��74�I��7N8�O<N��[|���>��'�y��W��[L�D��ۭ����l�]$� �9@HbD}�2|
��)S���Nܟ��<o�y��cʰ�X�~��W�l�w���n���+4;�k��܀�=d�V���,kA���-���N܏x@zl�6��B�˫��
�ߊK���������g��i�I=���зG�q��n���K���P�575��D]Y"�A+���,�)R�lj�����Z|�,M�N�|����]�魀���N�$ǌ0�7p#n,9�i�Ue�;t¨�3�ܐ*�Gp��q��HF��Wf�J�H�U׳��#�RmF~��4F3c�?B�iq#�[�p��hϔ�{%4�+<���C���Ӏ�婶� 63m��3���G���I.
o��q
$tu��^�ڳV4)�:9�J�M�z�\�d�f�I�˿�be�oi)2=Z�LqM�Z>$�d_/x�'��s#���	�� WKe�������p��feQB�� |��͛ae���&$@���q�>|��U�@~��h���pY��ѿx�A�č�n�]�4��Z��g2튶/3�'��m��y�����ڞ�H@�:W��H�8�-;X�͓jXc=�d�&	
�ΖO��[���Q��y�o�hm����Q �$̾P}g�Z�Gf21����'��G����J�4T@� �2@�_8���n'5��:��g8@9�T�-}]Q6�a�ú���9��!`���"�W%!����4%��8PrßR�r�p�(�&�T���')�+ޙ�u���Ra��7���D/1vm~��C�pF?�h�Ko�V"m����FI�QBC{_��f�B@p+�(��縗f� {��T^�[�7�R]�Ӻ�|!9P�:t���l<썥��"��'���@$K%��E�6�Ѵ_�L,��Z��b8ߏJ͏,�H��bx����������z��O�u��!��MoFC�A�<�*��-���-Q���!�!؄�^�$88����e�F�^������3;��2��"�j�#�h��n! -�6�����Ҙ<�T�&���U�_R��F�Q���I�n�7��Y: ������O�7@z���IP9�B���)�d���v�g��#�ݢ�2����3��g��a�?$KQ���+E&��Hv-��H6���2v�Z\a�����ˍ��ɝU�c}Y����G��%��BuW7��a�����#�B�ӟw���F	�x����i��x�46�Ok�:1[b�\|?���_�)e�2vy�C���v�_��.��~B&��J:�^���o�k�0H�3��Df1\���O���&֢r���s�v5����M�D(E�?���:��o�+B�`G��e��Uw+��R �����v��'�{�Lq�*�qm;ZS2�z�v�G��ޱ|I��i�k��h�/��"_�3�/��.�Ś0�W���h�T���r|��Q���;���D�����{6Jw�-4���S����¡��a�@g�SIؙMx�	����4� �^��Ӧ?EFl���4����V����s8_�SƑ:���7	!hty��]� �z$s2�>{��i��iK݇����'
=����~` Ȁ��;VIL F���V�-��ȿ���P������ˇ��W*s���X���A�>��p�R&׼��,��x���On�d��XPl���͵=꠺�;tKշ�fꞀgh̠Vh-�WЉ'���A�R!*��$���" q#�Ku9��Sb�2�Kc�0�h'�D�j��MG���h�0�
�pI��M@֝k�z��0�3Ҙ��<O��x:�����F�}bk�2;�%����a[��B�=���]`��r}�H�9�׭:s��Au�
�+j��wY��$�-�ftZWȳ�l�l�z"���A\�{m
}��C�&|w�Pv�V+t{\� �v�{x'</��I�bh�'��ۮ�q�����ա�D��w�m��J�8���L� ��ee�R���h�ݽ�Q;�M�0哺T4|�N���c��+�U4�b�,"�ZYJg�n���V��H��Nz�,��$�cx�W��zl���u��*4�c�����v^��� d.9�D���QqOχH�N��N��+rQ���n�����C�����\p�(��G� a������۞�3+h�$�ޱD�?�9���.#�5�����۞fKV,�����o[�U;wI��.���03�4���EE}pYѦ��ވ�Ҡ=������y{�6F9����D��3`��ZK��s���Nh!���k�Mȯ\�#ψ~��̊�:<�* ��e�_�_�@2Q��*%��lΑoS,�4��(55��_�e���P�=R�ϓ�0V�/�A�G�0aM�V]�}���vv�_Ǆ��X]�!�a;|�P�v+f ��*Se#��0��W(�ԟoTi&{<J�����%��2�m����_,Z�{�)��Q]��H�qA����#�4���C�<����`����3�P9��Sf��-2l��U1t��2Oխ��ئ����>�	\���i�1l,�-�G2� z:���K�b�(�g/�ͽ]e�k�V�o����߇�X�5[D*Ĕ�r3l^���ajሗ.2�}��k������*����}�a��]����DG�>A~�i �=��G�l;�s��,݌�\��	��{�d���{�6a��߁g��f�����:���@��6S\2�"c�QU��\�K�Cz����� Z�q\/��}P�R�{#�{�N�}b��\�;pxMN%�Z]U�;�MՔ=Mǵ�T�~�W*���4R�h�@��4Tp��eWC|�Z����̧.	Ե>I
�ys��9(�\��>$S���[t��l�}N�t�lD��1�p�⾖{�i'#b��D!��w��u�ڑ�ܢz����J�Of]i���'�5��.�7��t�1)$$�/���9\b,�Ю�<��R�ͷ�x���32�Ӥ�ě̈s�����3��/P!���Pڽ,,`j�Y����E�Y����ס��r}���3{�C�mz{� �����FQq�&�Bv�Lޚ^�v&jz�;bί��f��s�9�j|���9��j��-�k8��+ڟ'F3����Z�;��O��@�Y�l�8I:�4�`�-}h����(���s����M5�֓�;��UJ�Y�h��_��=�Ϋ��&��z�rɐ�ce�u�I�YO�3��o�p�����&}�&L%ת�ҥm��cL�,nF�� ��rJ�шG�e?}r��@����NL�P�V��}ݓ��U�%z�?�09�e`�]� ���ȿ���t����('k�c=��K�����9^j���O�'�L��v>�}\ڌn����h�y��ٿ$|�gCo�WW���3&�J<}w���߄]1���U>�����TTCe���Qf��C_��^�5�в��L���e��XD���#��c+����$��З���=�����m>d��~"���\lzQ���`����SC��ܕ0��-)��G^ooW�SN�}|�����Aq$�.4��o�'�������T��vy]�p4[n�����.�us��D�E_�C�G�<X���iV��<��C�U.!�@ٰ�7sj�w���)wؽ92�mPr��v��#�p>.Ƞ�snæ<h<�_}�kʂ$W˿��2�!h~����IR>�}�2�$���drа����6xs��Kx�믁�;˟a����2=���%���.N(Z7�7K^��I��RV��A��8XF�����;�:�$9*�宷�x�iqtG����뮛�)��*)��{u�e�9!���!���45�ﾎo��H���bN$n����4�Y���q0�v���A�Z��ס��&J֤�[.��x���V�ߠ�gȮ=ݭ���m@���{H��,+8VX뒞������2I\=dZ�C�.-��giY�<x�W�T{���9�3�*Z��܎om�ѧh]��:�"��;��l�ə��\^��؏}{O!�p����*�y��VQđ�L�����s��t�m�̎s��1q�>GM�+y����F����_847�آN�HR�%���F����D%B�Kd;��2�����`خ���fbe�JY@�q�toL�|��	��j�����p�J�G����o�#d�u���Q���^3Z�@��Ϝ��U\��ncgș�!=p'�@��˂�=1�D� �qK�\���)�@g+͞���;�I�*p���X	?��#Q���f�m2(r��4�|�'�DT�y/����AIթ,��xX�f�`�0��� As�jd0p�H[�cPިe@����Ĥ.���5Ѐ�y
�X`�n�w��*��w8Q��v�^�F�M@���]��R��
���;;]i�E1]��K�n�ȇ���sX�^>oS��5+�]��ӝ�s�
�w4�x�6G��l6楦`�|�[	��V��s3��C�Wj��A��^�=ً���[P@6��Z�1si���ېk_��Am�����65M��6��	�J}ͺĊ���>_|�sL���o{�5��a��,N+�+�^�t��.dj��-���%�C���d�9����Q�F��?�,��/��-�+ۻ�{G{i�"F�J� =��"��і�<����0|A���r���7m��;\>5��l9
]z��&g��7?I��$����JK�s�����.�����it=��F��޽w��{�M.��� �̏;��$ͼ҂O0W�����pE-��2"m�����l \�ں��JW�3�l���هga�8�aE.~������XQ�#�V�Y�v��.,�6^�֕d��)�b�<u>H�,}۝�xf�TY��+��T{7�.��2Y�mw��oy� u>��tjyѫ������tM��#��&���wK0u5�d�D��<_��T2��l�}b���6��]�b���3wl�?��&���m����Q�Ha<��5zHrrv28亡�:|)�
$��:)2ć��t�ŅY	U��G$`�R��c��k�?S黆�RlW��g=��W��fӓ��dҾJ3�Ȝ��͇����L�ȓ��T󋈣��YR���Ǭ�K��F�C%dOS��a�e>QH�8.�|*�uN;*~hD��K��y�+����t�v�^��U{�l}{l���f%�MŅ�*{���c���U�ߊLn�Nz��)���y��#�1����:Ol�nI�Lm��3�G�"
,�i����=\�S�x{u��cJ�b('�q�Y��ug���V&6��1��y�!~�t�o��2����'��z4ݘa�+����\���	��J�vu�1��Nyɨ�xl�If�\�ע��KS�
D"�j;��c��}o�"��C˙�����/{�x���~f�'Mu����L�N�$X��iU"�k6q�in�����d��B�dt������PZp8qߐ�`�+�1R��L��RD��qj����&<����}������nh`eկ!��u�z�
daeW��	-�������(>{":*�ֺ�ʦx������,^	6���~ɴ�'}��	�����I�r�;��p%d#V����/<k�8�W�]Ȑɇ���Ϧe�Ad0%�f�Y ��D������c�*���w:�J�ߤ�*k��{Y-]X0H[�k������x��{�J-
��m�O5^,�:b�M�N�W�����Xi�Y��\����w�K�1� ���ɘ�~RǞ�г�C�\S#��uhE��7�d��F�γ-�b�zHD��[��&,��	�&k9|���N�:��n�cռ?�[�;�  �G��u G՚F>�V'�53�,^`9uR�-�\k@G]�3��Vvamhv�j�w?w�c�av!]B����0��ǚp��O0m������=�4���6���}�|����.�+�tl���z_<uР"�JL�/%���O�]������������xJʱ�����/�A!`�I~�c��0�� )��?��g:��AUV�)b���](���JtK��|xF�iu���|��i�+K�{�K��z�v>|9&(�y�Mw��F3�r椷S�6�fӃ^
=���]��AH�=�]�w��^������ٙ�#?�;��R�ΛWs�-��Z��X��.�e��4	Z���KX5ׁ\f�0�P�'��o�wp.�+��)��p�H�OqZ�ܞ^��o��S����7���})[)�� 띦�՜��u�:��.W�5�㢾���C���Xn?s	J�������d�fއN�Oz�́ۉƈ�6:α�V���c��t�8A|�&:;��^(�䛩8{-˱�X�x|i}�qs.���`~�t	/P�C�ޠ�*kll�&�K���IrY��_��V�*����,�gC*?;|;��$��\[9��g����%w�-3rf��RS�����\����nwWh `�����<jqјzg�;���Z<��3�Bu0�C�=9�.F�#�4����p���۸
�Szj�O���giD���AJ��z���q.;������
��:Vg��T,1�S���e<3c�97W����5�y_w��S¨F�G��c��bC�۱y|un�O�3�/gؘ!���8�A:E����崴�-9�p��-�C��"��;�ɧ�+r�b�O���&ú�E	,�o�	u �z�S�E �'~�n���u0g'���e��Dا�Q��w��a�)7��� rX~&�Ь�?�;�����4�x6���>�It��^�h8�z�RK�y��]�r �vF9�.�%}F1�IL�L���ћ|�_(��\E+v%� V�/���EF{�^AЮ�+wcm�|�~���5����3�V�sl���q�pcJ�).�b��Z�sK$�D�9=� ����U܊�N!K�D��?�������^B/ul+k�o�t�>����c�Y��͒fӗ����������k>�����˱��6�rR�ih�T<���+���T�o�Y;?�tF0XC:��xPC��R���gjs2��e�6�ɒۺ^o|��<��ڻ6ј��L:6����!��X�x~���5L�Ce��V*�m�'����1�nl��;�T"�����LZ�V�H��GQ��<�Ψ�����!��@#4&�r���y	������{'b'�f4rJkн@!�l�Iv  �+v�u�c������2.Jo���iD��k�9Bf�"�CR?rCՁ���n	;�E�Oy�үcz���w���!��z�։!��7�A3F�������y��K��x��l��;�ʐ���"��;��;��r�����~��Ր��f���d|���K[&�Уry�!����^���H�t��2K=I�=���G2wD�e��gg�e�;�G�-]���q��?1��X�����=��%��,9b^Y���9XE2kS?���#��������xI!����	�z��e=��TN�O�*��i@��)��U��c�a�����.&X��%6���æH�[7��V�dn.��U �8	�f	|=���Ϲ��ƪ��gGK���o5�ͫ�}����l�=�U�G�})���f3��k����p����OϾ��L)ra����묁�� ���� b*Ӿ��e�[M>�3�!�aGҤ�JH�#��چ��}�V�ڠ6���#M4��\xAXi�y�����V�*ȭ򘡬���� ʚz��XD��y����S��Vs�4�j��� h�~� w��Ք+c��b��2�����+�_eW,�ښ�g���B<k�^a��?;���3D�k*S���}.G>M��$D�����p�F$`~?;3 `��Y@�7\�[U��^���h�+<�����?��jR(ͦ�x�����	U�Ϙ�\���KM-$�^�o�Z	s	=7�bj/�;��>�k�͕�G�l*�U�r�#0�8�q1T8W���﫩3�xݞq�6��o~`��R%�t�3ᖄ�q�Q8�:����		�,�Z�L�&�����5��?�O��Á���=���WR,�p���be��tX���j g��K�\�U,�#,�f��s��Ba�%���vM�n��ڔTL�I��l*����!9�����P��и}-��8�~��
#��̺�#������sT��ʕM��%��8��NI7�D�����5"��v�coӘ4Xp��7Ph���5/�� �ć���2D(wW�2v[�KX��'�R�x|nm����7JF��)����s����|�y����>F�v��)���uc�klx���z!�Dl7��%-�Uͬe����v��yl��_��b�!TJ|T��.�E��M!b�S���rWO��+7�[�X�~&u�-n���q��6=�4h�<����Z�J��#2�'�	/m���B���oI�Ղ��G�b�����P�I6-�<L�}�*�)�f�@��ɝq`��ƀ��pb��i�աnV�7�f�,�$[��^��j�~@���^�0�#UYqB%X]M�����<ƨt!9�_q���'qrY$�����h���6��<Z�Z~!��e�!�� U���� ��Z��q_�5�{�Z�Hp�3�Y򀩒E�٨o�VGP���8P���[�J[>Mό�hy>i!tcsq��e û�o�iI���IG�n��R����C�U�p��&�*��襤�5^1v*���~vVy@$���/�4
9cT�uP��E��`�Zn%wQZ�B�X�N���ݘn�yX�|�������!�G�~�Ϥ�J�v����ٖ���ia�����E�%<�s�����~��3O�ҙ�v�V;����@�c���+�*�;M�nQV�	W ��5</�C�{�+��sI��V�s������C�S��j�>����T�w�v��f�L[OM���l�lt�*7˧��|���B=�p��}K�{�@�\Q��3��K^vr��|�p�[B".�����*��iU�شp,����%}�&g�N�9�U$����ݿ��z�+*(ڽ?L	G�<� 8��k�6��Su��I'���v��nO��{��YTԚ~D8��~�v�J��˾�������<��[S��iP �r�Q(����I�n!�:1C����V3�`ھ���R���F$����BMണ-����ĩ�;7#�χ�W]�JfM;���يf9��K��/a5�@��6��0	dLE�)M�O���囘Ҡ;�%���d�L�}ir5@�*ܦ^|�78wV���>�>�T����}���g=8Y?���B� �h����v>؆��9���
t���������V�3a![��1f������X�6..�A��J?��D�D�fP�Lw�价������{�u��%���dX�	�[�����Ý)�د-��e�{�ꄄ��b3I(�c7����+��n������a��-O��V���З���+���a���"	�L�@Oo��m!�]�o�^��n�V������E�rZ�UN�F��#N������ύ���CRa���)#]�����˙���=b�����۱��T��Mk���{萺:6�"B=�\��z��@�-1)I��%��|�����z��k��ge��q��qҵ�Gb�{KwW�y���6�qxz�I�I_���k:�tv��N�8U ��N�QլJ>y�z������e���pm|3�ZM��0�S���G�%8�����~a��G�Kv��):TS4<�	p�v�t�1�,�_�-���||�Oq�h{�ϛ�oԯm/�1K5�C6��)��!�Xh@�nT�?�=��_>��i�br��V �_��Yu�A�F�lOSs~��J]�|�ⓁdIm���"[ev�ߞm9�<��gO�S2U��5���KG�7 +	1%�R(���B]��~�-��S�<��G����t
�+$
��b�c\����ռR���AK�̈́n*�󮱵K�H|�Q�Y�s졹�.?�n� �R9��*�Oe9�N_��oB��?����B�Gf��x�'��w�~e$.��Ưlb��7��	^B��
J!�g��.L\xA�2ojatA��%��ʌ�\����i�I��������a`L�yNVtȘj�h��74Lc�O\ nA h�K��x�J��Ç� �D9��V�l'���Q�:�z{�U&�?3:q��W�?,0fA���M�����2�WQ@ֵmtgL6�`Cᮔ�(��� N�H��:�e�4T4�>n����>��F����[�P�A"��N���|�'���2�����wH���ϟ;1����Ӯ�ۛ���Y�g3y������I�� � Q=�[�gHstk��\93V�^s��T$���n�ɘ����
����%($T�#�(FW��F��r����T�-a8]Rs�ӻR:l{kވT�U�l�I�8k�M~ʞ* �~�dn�]��m�O�w�h����gtV��
l�ig]ñ&|��IK,���dM� ��}F����@�UP*ؔ������Sjj���rN���N�d�T��pW�O����*�5��c�â����QDP@JAR	�F��Α����D���ib�!��$��;��<�������>g����^{o�K�/ ��p�n�&#��;�V]w�����n�T�n��S��7�M�J�H5������նGo.1Z���?�C����~9_�:�TM-�d�H��$�m}�[J��
�z�Id�L��h��ni\s��d露 �m�.&��8Q�>��7����h�ꃜmY���C�����ӏ{xU��)Ȳ�I{E�󉽺��L�� QL�XwWn���F-�\�o�4K����2c��Z�5�i�,�T�kڳXJ1��F�C�[�&��C����֛��+�
�	��y}%�<t����k�R\\�^&b�0�v9�p��^� _��̒��KXf�[��a�.w�5k܎%O+y//�l�;�m�޵�"�U���W�FtJ)\��3��I��R �,	f���i��mޏ5��z)���t�Ҿ�����"&l�z�:5�\�(*�`�W�F����T?�SQx��Ӿyg@T��t�<.�l�dw�6I�+��:J'�۫�S�V�#����t����Ώ\�݁�o���&m�h����ó큣o��ioI^8"ޠ�q���#erfhRV�[K7u�v�H	�&��7a��j���lMJ~������y��̾�o=%A��q�]�^%�*�> �65=wy����SX|�f��=M/Î�-՜�@Hǟ�S�����ѣh���+�~&�g��~a����L�l'�����Z�L;�I�M54w���f���W�u<�Ϧ�t���pG�DW��o\x?�B�bO|��^J$����t}��4D���d�~�[�D�O����M�+��ۺr U��T���B-3���؎퇣g����۸�j����,`~��*�a�C�W����}���M�C �e��E��Tu��q~���W��v�A�I/̫P4���x���u�[o��K'��d�mC�����[X�NKb��V�_]�r��F��Q���1��cY�����Z4��8�/'��8�0����-Ѫ=DgMX��s������Pw��)@��"�Ï�؆�O��Ɔ*U958'[��o1�7*s�rbп�/��ر����Ľ#⟬8ԍ"ӝ:�_�����h$�u���ER������Z��^:'��}Ӟ��~�������[�7MI������y��n�����e��;r��F[����D+9ܓZ�FW+�b���^V�ֱ���|�8���>�z�k.�:΢�b��2�0i�;���H.�'�
-'v�N�j��Ή!�W��dw�����1�w|��-�����D%r�o���dp��_�'9�'�����"�M',8~iZ�,N�FQ-��w ��h�� �0X+�
ƥc���)�^$��N��l2���߸�������Jg�H-�9��#��i���~_�F����f������e	Q��v�ʭ�mh�r�5�3���EC���{�a�gktk��=�-�����L݂�`	�[5m���t�'e1�����l�F�*b������dJ���a�=-��M�Z}��2r輰��|�nw�Y�py���&>}��x�m��%����Al�B��z�O���t�L�B����i�nOm�Ƴx)��o@<BZ�3l�g�K�����W�򎄋O���G���� Q��5�਱C^����X?@���΅&�	�j�-"��C�m���t�FI�
�ĪK�͵�$ej������F����)��<U&��^�%SL�$��\�=���^֠�D�-�]�Xţ"-m���3��S�bه���G�8Ḽ�S�r����lި?;:b��7�.ǔz���3ti۔��?��=P7�}&n"�{fjPk�ݢ�\�E�v-i{�r�G�I��	���W��-�c�Ddp���^{�R�&]u���ˎ�K�!#<��Hɑ�-Ȓ�Ї�WuI�5��~z�f)ξ���� ȵ��n��I�/�/�K%'�ҕ%R�O-���a�+o���ŋ�h�ܱ��o~!���R�r(����h�y�S�{��b�P��+	f��Dv o��c��OW�qv�Ep\��[g�j���+�EF>���}��*��n�5�ۧwg���rw�>C:�VG�w']�F�ւ8Լ���� ��y張%���cn�2��F���@NA[�w"N5f҄_ԶT��,Mz{G2�-[���9�m^_l7z�{��.Q����g�+��̭��y�nL��Vх3��֧�9@���d0Mi�w��3��$گ�LH�d+Kˁ4L�g_J�}�4�˭pM�
����e緧�dBX\hr���u��"� ��Px�[j����6�R�7K@�2z��ܐ�l���Aa߳WEפyM��||����s��y��,�`.���H`�a;���&?R͸tOa�!,���6,�6�8�L�{�;�K�����o����U��c��$SY��}O���˩`�AR�{�������q15��W�H�J�Y�)j8Ơif	�ʅ�	�b>x�Y�P}T��֠CrG�Ϛu��~����qLx�,���
��}����v�j`�`Ũ[��G��qQ�ب`z��uӄ8����{e�@�K��]�.���M�����mvw�T8��SDJ=�I���xϷ�o�;����}�.4�|d�R�|�#L�:ܞ�(r�[�� �V$���g[���� �d�̽�W��d7@���4N~�|��&Цg6�A2PC6��� �q=#���E��� ����8��7��,Iz�>����q��X�t����/�T�1����I��Zf1�s�/�~����d�:���4���a�h�Sy�����Iyw�Mx}�U)Mf��Y�ԥ�?쭣�N�˕N#��v�/<Zo
����LoDtQ�p���X�QC|���ŷ�H�rJM~��#�;ـ}H�fJ��M�6����:&7þ���&���!(�n���������U��CR����h�O(-�r`���o��c�V�����D�өF��%�D�ʈl���n�s
cA	��6��8��:8�F�ܯ0�߱�q��!!�'-�wah�c��J��j��VV5�D᳐s���K��#A���=E��7��̻�7���-�$-��<;��w">�t�s'�	�q9����|��ӭ!�-���\c�']U��eG�pPs��\72�����N�P��I�v�����m$��k�|�_��G�T���TD*��*ؽ�0��T�JY_Zx�����:���j�L7��(�scaQ��k9Osvq!'����;<����.�m��fa
K�����)���C1B-���	ub|�p)X�hC��9Ŀ�r�8��`�j/g�����ظ\���s�Ol4������E����
��=��2��E8�Y:�cU8�&(�LK<�9���n7n�uç��X6�� �/�z����I=�`D�?/�]R�AOH+�օ!JyCe~�@���U�/0�Jd8p�Kg<<���Ϗݷ��ĽV"�>��J����&�L��Aiâ�gK���Oy{-I�	�w**��%i8��r_��Ⱦ8���K������tk)JGz�%:��۬C^�2��(h�U��kLh,��eY���ي0� �~��8\�dW�/Z��%���^s���~=,��(G����VUJ#{.�n�#;HZ���,�mt�	Δ�}q�I����3�@@�������}���Z�E wk^���2�H{��]W�6��iy�O�9��p���oZ)��-��ǵfP?�<n�տ]�$s#�Ȯ��q0�(�u�'�|����щz	x�j�)��x�x��S�?vj ������{d�Q��Sd�c6��x@_��Mg�	E�TZ%�~EeO��/d ���s�l@6fLa��������P̹G`�5����+l�B��0�/�B�߫1�VC\�ȸJe5|���)��faҲ�9a�S��\�*��F�JUW�e����9N�����$x�ӌ���%U��c��
��0�Y�����y&#���X�=['Bt��H'�-jf��4zI���f[�W[)���������U~�Y5�Fn�����#w)��C�B�Q���A3�h�|?8�%������ݽaӐ�K�?t�&Z��G�&�4W<����g�}a���@u� B�]EcjLC�C����H�D�R�+n��{�\���:E��9�m嬥&��!�Z��<�[u�{����$��}�Z�
�P��a�K�%��Z^�*��\V��/,`������z{ �����=����n�j����=�)�%�M��Vur�z1Kәrq��Y�OxĵR�!|7�'�� ց7�".~��T���-�$�;{�ȣ:d�`5z��h��MP��_�g��"$�U�X�S/�n�=^��j��j%�/��o�c�v�뼸4Nƒ)+=�E�A=��ba��|H��BM�Z�e�53d��S>�\ż���S�^�9Sw���#7��=%�F�<Q<aoۗ0�[2d@�M�$$4v"ė���k��R P�tϟ��ꁸ$_Z7��i���^h�k�nX�����I�I]������Ȼ��ֈ�ɰ_�;Y6��n�ʻ3����	\n����������1�\�e�Jq~���jB+�D���"{��
W���J��s��/������W�qBGme�Q��7W���u�Dp������p�Zf�P�N@y��3GY��A.q��T��q�%�����BM�]��j��ϫ�,�Y�F9�~v�y��l:4�M�t�b��_�=�(%������}`�������(�����T��q��2����G/��1��Wn��L'���jz�_�b�(9��3���/hH��q+�;Qx$J��O�&,\���Q��Ҩa��>����v��̢ח�s�:D��}D�x����.B%����l�Q}C{ ��d��C9����7A���K��8�)�z|
��)��d6�ۈ4�s��r���Y��ဓ�23����
9�3� b/��ǅ�1���l(��A�7�����L�F����k��z;��/Gg�x̣��?cbW��r���,zEkz��I��px/��]�5�$zM�F%� ����s�A���2���ez}ݜX{m��K(\���?�0�'�}�f.29��.\8��U�\=c4ut�T�c�0j��x����X��U��
��=�AT�@���c���[��"ݬ��M�0T�4b���]I^�K�nS�?�0���cN���a4V\ӏkT��UŖ�oЂ��㷍����,�����S��=ψ�r�N/#9'����3Z����d5�I��
���W���[?��PXC{�:r,a�R����"�Na3yQum�{�b�\�)�B�x9�z,=7�T7�KNp�JDbb��b�x�洰�����vD�#���B�V�8�6�À��[a� I�kq����;k�gQ���ۏىhO���;��:��ɨĿ�S+��`àQ@*�ߚ�EtǗF���n����{L�AD���[a��"�o	O[�/ �o�9����	��A�f����d���+?#_t��fqn������g�Ʊ٬%9O$��*�u���[-L�*]� �d�H��"!b��3�C��먿zZ�ڮ �3�V׼Jţ11/?.jjD���B�z����=
�4+*rn(4Ϸ�d6�7�����K`+u���������F��&pw-3�;R�f��i�H���瘠[hb�@�q��G�&�:�_:�� 
�{��(XQ7=L��<&�m3È=UԙQ�DY(#��CZ?�ƛ��Q�I���]w��A��g]A&���_y���;"P���)�N:6쟫�$g�S�,*'��f"Ӎ���l���sԩy��̪)n�{k3�2�-���x6��B����Jn:
��k�55/�R��0@8���ۨH��/KT����>d��ցd� \�@?��n�o��V�'
x�Tg�5J�M�<N�QAw�\\�De���=�N'VM~�A梪C����a�c�@x.�##�w�9U@/}���j6�q������Q���o:�n����ϕ3Jh(TѰإ��U�C�W��n7�/�Iٽ��M-3B�(�?��O�R~,O+Q g�����ǺĪ�j.BH�/x��x	�(����k �����ez�Ż�q�Vl.���K������-f���̰�k�:�Đ���� @#q�/`(�РRL;q�ϳӚ���
�_\2�����ql�B�:	�:�d���y�G�U����H�C4����ʸ3�4��ޗ��7f���<�T���r�Qj0@�����6((����Z����h�3J�i�Uv�6c3;O�Q��ɒq�h�<!�ʿ�:�G�i��M�����u�W6:d�Y�D�:���"�)���TCkh Uf��)�"XpE0z�q,�lѓ�J� ��`�Jퟨۿ���L
 �1��w��eg���#nf���J~�H���5*G����i6"d�}B������
3U���K����6��,'7Ξ�F�������rO�����?!Ψ�N&���k�-�U6�<��h�O_W,�0~EŽeE^_{��C*i��A�`�Iw������z1G�>$wjQ
6����g���@�}p)y�{�5������k�A���{@���?����d��`��۾jf���{�A�V� `<��2^�r�Jλְcf {�v⿿?y�Qs�'x�}5�Zd��sv>�=+��uG����Z��p����� ���ì�	�s�{'I	�le$���/Dgss�"2*WO32�/���y�l*�lIX��a_o|<���I-SG�K9_���Te�l�](C�a�l���v�lآ,s	�~U�=_%� = � ���uӾ���Ռ��f�$Ѵ��#C-^��"�p0�*��X�Y<�LK6���v|r���ĸE���y�}���%�t� �a��l������0`P�d(���O��q�)o��t"�<�q:����A2 @Otl����ChG%�&���=����:���VI��}����|4���৭Swf���R�(�-�T&O%.�z��쏩�
B���� �~i��0�>����	� h����N�N��Q�&8+H*j �!Q� �^�� Ӝz�j ���\�5�rQ��'!��7A�'.C�{L=�.\������ ��K�Jw�aR*��ڍ�-�<�!S~깚<D���a��O�� �p�-�a]���g�L+�G�wq9�%���߲!z���ZX��sjX0x�A��B`$0Z���`&�R�p��e������c/̆K#���gL�m�ŇUh��\���s�ل�S/���x
h�R|�T9�9�~ݔ1k�p��D��OU�����m�A��m��e���G���w������0+�z�ߠ����O��Fr�����5w�t����\��W�D����[��@|���JU��:<{�O5��墎~Ң��~z�o-|"�@��D�z�{�@��X���u3���&1 �@���L�H]�ss������	Q�v9{Vx�f���;4qh��Xb�� 8ė��G�'QA�4Y���B\�B˱H�},*�\�?�b�v�� �ӻ���c��w�6��4���H�s7����_���s����� �x�0�Q?5t�#;����X�,p��q9/w ��$�Yp���:���7�M>?᧏�������&�mq��h���K�Lm�/;?O���-;��,��c֯R��[W�)�� �+��4 �䀦D�B�9;b���)�w���oQ�ZP_��� b-9���p:����r�Q��\z3�N����r��t9n�q�����q�@/-��J8��9��U�^G���5}tGt��i� �ϳ��&��������;k^ir�$;G�ql�^������Ա��϶��(�h�f�!'6H��� �0�o�%��/G2���r��쥓@|�8:�KVSS�Xdt8;6�.���f�M���f����#��^��{�a�������.��X�?�cz���CyrpT��>�{�K9: ���kArQz�����"2A,�|�;W@���7�`&�)�>^����9.H��d���v\l[]^V��i��@� &
-yӿS�-hי����R�'3B@?���m���kU��0&�X���h�BN�1O; ��B��"2�2/�l���z����H�O�z��0a�i2�7_3d��Ц�B�w�2�2��Zeӄ������C	E�
��^����~s�'�l"�t����F�m����$ZQ�����"�r�F�k.=��<y���Ta�|g�^�ċ��銶��q�W8�=�P ���Dk7�Ϝf��z��V���)���i�]7�O�s[�]�r X|@����D�o�	`ܤ��8�ߥ ���������n����sv@ԧ'��j	����皵��d�����{�:M��|/%�6�O�M�b������7�m���܉�%_ڟ�6��-A<u�^�v-f���Н)̲[��~�P�������#���Ωaӄn(�ڽ��%cO(��b�����w�s\�0��9)�i����[�=������	��!읃:#Rn��ƽT���$�h��K���VbJnx��4�n�9��[]x��I 翽08ts�}e��O{)�%L�#W���o�R�o�D᫏O��HG��;/�8>�J�e�1��[�h
fҤ�:��Q�6m�����y��J���N���}��2r�#�ź;)B�/�£�����U,��͏Ҭ���A�����}��Rx��P;���٬i_���.7>���qM�z�0�ۣ��6�؝�x��(�|'n�\p��+�
��| ��S�Jm����Em֎�dg�g�E*���i�v��S�tM������������TQ%`ذ^/�--�^-�0j�qSD��Ɛ��]���F�/���K{yy�p#Xg�'s�U!S�`���	����qs�W���|�c9gꕡ<pf��ڱ�<{-��|�s1�9V<u/��{��݃K�TE��e:1Ҭ3�����É�����ł�o6D�����Π�����rb�͇�-����#`�>Y*�:�����v���{����Qk:81.�G�)dI��&�������U=��!H����J*�,Ü�Z�d��U�]tGn�`�qu�K�~:^3(�iK��hy%�?Z�%�����t��8Ё��/�(���Q�*6�,�u��1�m}-r�C1��y�|�X�\��k��HK���ޭe�{��.E��B��䗛�J�5���I�`M��
�z���j��YCi������>#��
1�u�H�@k�TWjfc!d ^���2�6���]���",��#0/4��KR�	~���fӽ���dcj��%�J>$����(oz�R���$}�U ;_�r�ޛ*t#^�<�ՂLik��3���S&�E�%�:��X̼��w>ꜰ��>A��B�恛t�3�~ᠹ�I�g�`,N�	+1�B��;�i�T�C��6/9*M�`�b�OL��� �z/o�?!�)�:�q�EY��Ch���\���4���F�@*9<�x9��@�����n���ݞ��ڳ�Q�"��.�j}�- �&�>�����cPg��s2��nH���M3�~l<�������\�::�"#�*��IH��������q�WᲑl���~���"��e��ly��+�$��g�nOҖܐ��~=�q�	Mѭ¾*۳�%�\lӭ>(��-��ĸf^]*���wŦA�u�lb�1�$�U�M�"ϻB
�LHDӷ����KQ��:�8�~��R�/E���m���r��.3<�Z�w�o��~7�(��v�C�5L�=	�^i�G�HdK��,s���������w���A�"��O_`���՜ ��n��j׸���&o�>��0�%t���vUS�s1���ɆM��Ns�[Oas�Jd�8�������l;'v
e�������6�<x����α��rO|�Ǿ�}	��W/oMߪ�qB�
���)l�SE8S0@�*k�����!4��ߚ��/�
bk�>���/	�����
S~Bq+QΏ�kE,�~���x�b�f�M|!���e並}�g����uS�Fop�N��T{oT����-`A��(�"lvFnT�0�؟�w�}}K��
���h�]�̽�׎1W/;<E��Vⵖ�t۹E؄�����)�E�&f�Pg�����[��zN�~1�q�b.��"j������?SX%f7����.���N��m�W({�^ܕYgCkP/B(?�J#�3<uB���&��E�ر���̔��,�nՙ�z~��K~F[����;�Ćy@���������� �K�hBn��s��=e�{FB$���l�x������B�,�%0( d�z�I�������(��n�(�,�ƹ���[Se�V�^l�k'^|[oӵuR��8��6�1u��]���(�(�o���c5H�=E���i�k;�G�����hX(��7c�X@_���Y�($����u�#OA��[�� �����+E�n\�A�Y���{|C�'�����%���O��NLM̨��C�d>���hS��4= �X��E����gr��IU�,8�������ոK���h%	Wo�%����j��Y}5�l�ҶU��>v�7�e�.C�J#9�F���R��j�������!�8v��CW9�kW-�%� �>{�b&q��#%�I[��6�uq�e;tLj��,�����m�·N�~��=^�
4o����X�hJ��Q�6z󚝪�FxĴ�p��
,�٧��t�F{�o�.K��b�T�Z��K��l��*D9�:�K���.AdQ�w������ ��H!M�C�<Ϥ���d(��+��>�^Bn8 z�_M��n�\�t�dp��!���)��qa�8��Q�]�a]4SV{} c�9<���*�X�j�����$�tp)L믅/�����^ h
�Nɟ����C*�u�X�Ĝ���{u�
o��;��5T��[��ҏ��4V�
2j2䪑	��eF^:�~�.�?�s�x0��=��௪�Kq	�H��(;:y��h첋E؈E?E�=����Ƿτ�ƫ�.65�	����\��Ĝ�y6��6�O;M�u-��ع�K)�b��u����g��U~7Fz�[�W"��z��5��|��\���#��2�������Ї�x
��6m)�����z���Z�O���,q��g���FP��iy��%
jګ�.�My��7����b��k�/�ٗ�Z��65g��xe�t��ce޹y7�j7�p�H�^�@�TE�ի���<��@���֠:��r�V�^m7`��*j��%�_%.O ��7QU�+T]�r@�IT�A��SH�MI}7Y������LY)&�!k�,���W2Qa�U�0�ח(R�8���*M=�ч�Wȣ��NZ�<W��#�b���)]� J�����`����z3�WϠ�����]����d���x��G����*jF�6fgU$#Pd_DΛ��%��J�`��L��Dm����~�����z����b����ߜ�R��z�駋Ҥ�K����xصǼ��������ݣ�R�Fj�NWغ�r�uu^��p�=��_ٞ�7;�/�*1_�<�8<��{�0Tѩ��;Z���<�p���K�����q��r	������Ӑ^�YA�<%
���ң�I�K1�����aw�w����۝�+qPz���f�
k��i���Nj���=�)�-����(����B�{rÖ+a�p���%ቻ�&>r����U�l|��r
�y�*U����bN��T�'�bi�%Fi��Dl`����gowA~i���$��QG�͵_��r�Ʉ�2�dj��H�{��VXI�,��N�6�u-'��0����4���SXEe�X��R�m�\]sZq%����R�,?��𕙖;�[�7`R9�������h� w�L�m""}�mu��I.g��FߨhQ��rbP�����}%|a��9���H��q�c�D�U�n��M�>L����Q|���ܥ��D�vMc��#7�9�ر�Jg�ǋ�&��~����)G~�O��<�\����T���0jz���9��eӺ�s5i(H��������m�;��7Y��d���إP�8S�;9e�7O�{>�d2T�SP���{Y��>��~��c�{C3aoN��x?J�Q}�pJ#a0Y��Ļq�h���������+�3�`����T��9�݂z�{s��=��ݕ���ν:����~�S�,�Sg_�6��W��.���o�&ANL��Og�WË��YIoOlPT;ΝN�+�N������6���,���V�Uk$;l�Kc��A`&��B)f"�;��_6�s ��/�>Y01!!fb�^���T��o���r������~�kL���t��Oh2��jM�	�	��Tv��{�|C��};��U��]i�CZ��2-Y�ЊT}̴r'�>P��K�� 7Ks�3�ۻ�z�\*&o�vn���(�H�#!��+��C�ƥ���yX-�!�_�e0#���F�2-�jEg�TR>����\B�S0,3�Y�%�.jr�4�����3�/ߍ��:��Ys��s�}�H7gi������4� �^m�;ݦ�",�ư�xd�s������[�̀Rx�� l��� ��`\�n�aK��Si��N��)�V����V<���o'��v��<�l%M��!e?���)sΎ1��4�o�Dp���"k9եlɿD�bL�� X�,1�~	��/��u�;t���(�H����7��Lw.�������y���18YhTŠyA}�9��7����)�;t�!�K�$3ˉD�;���(*ݚ_q
;��6'd��Z�l�Nˉ2Y���}�i�����Z~����K�
�8Kq;�(��E~v�=���Nx
�/ߝ�����7)xރeV@���) c���S����g���iyt�)�k���PǗ��gd%����GIK+`%d;o%WD@5���N�b���7�7��Z��w\��T���O��P��f�붰��M�d%Ak׃f�Ղ�������n�b
#ʣ������&�����#� ����9V��2��/܆Z������;�#���r��F����%��-��^{Xx�1D����:$����Bl�
Mi��N��i:p��SL��?L9���S]� �40`n8}�I��ס�bz*��Г�t�q��r(r],�_��i�*nn�],������M%̓�����4���T2B5ۋy���0��Pn��xKôzK35/|�k��	58�Y��&Ll���t=�X���ae+��ث�չ�-@v�~� ��D۩S��P�/? $�/}o������p�u��+땹��D��2�h�C��zb����c����m���nn�����3��q�IF�Bc���ʽ��2>��0ެL��WY5 ���(K&��c�`������v�m0:�i�`�7_Z��������e�t��Tqp|Z8U�Ʊ�b��=٤�δC0�TCW�NFK{wL�k���zțVq���F�%�O�s�H�/���?s*�;�a�m��;-b����7�-
�>�J [6Ј�k�#ܶ@��M���T�*����x�2Zwo�y>��S)��k ��59��u߸4�Wة��.`�u�2c���p3B8�w��j������zy���/��2��j�O�I�T�/A�E�e����f)����^ d�
M��	�1	�U�����g���]|�����	Q�����8�"���������V��p��r �ma_�ի�u)
n<�U�i��>����y�ST������-OQ�ǟ�FĀ�����o�ޱ/z���*�|���,��R~=�*]%)���7��`ms;���]�hUخt]Z�p��~
ݪ��L>�S$7J ��m�.��ꧩ�?��_~}��3��Gm�LT�*�����9�m j2��3�]{�ZNɭ������p9oD���x"M�C�*�1��\��N���������Ti�R��p����')+!�O5n���#�h����:��q�!W\�0Fj��M�>(ox8�m1�>C�!|�ޕ��$i���b��k����5�jH��$S�C���\��C° �%�) ��5��S�4�R�\�IF�W3Er_	�{<������Wai�����D�q�X?��s]8g��vr��a˗jT�up���S{		+O��J��Om�6���������/;^�Yg�o�2����&�z����%���(�P[�i�4T�N�t"��5"��P��k#���յu�א��}YW�R�.Ԛk�]��V��3?6lS��ymN$�:��S���S32�)1f��ĖY�Le�|�"����$��
*���n�����Ig�3���[��L���s�(�#��1��R|Dҋ�KM�8�&��hKـ/j�P�n-;���P����@ˉOo��x��;��s���u���D���iK�|�_Z&>�n��!"U�/!Zp�̡^R������n��EGB诳~#�t�ۼ�ڞ���3
��)Ӟ'��f��y�u(�J�s�7�b�W�|uʾMx!��spl��+�ow ����D䖯�$"�@(�]�Ԫ�y�����)+��V����k��G��V��[�>�O�x~�7l�f �x���6d��ַ��Oqͦ� B�M9�A�&�F�U��V@���Smw@��uF�$�[�QE�m����d����S��3M�C@����A$�YW{-c����R�4�S������b��>EB���9g�%�;�"b ��m>^K'��B{9Sތ�r,�����d�0?)��Q�������XIp�B|} ��ޝ��t�D�bC�O.�~B6Hb8��C�&=��F^Nt.���Ꮗ�L�˻�\�=�S��ʫ_�c�����v�J���0 ��u8���s� J���;V���
�+Hx��'�/���u����a[�dr�
q8�#�$�f�C���#MB
~��:;�'�&�����A�i��pջ����C=�=���;�.A������9�z��r$u-W��Ia[2�h���x�-.�V/WYX�H!���A�@x��Q�HE"вQ0pe�~�J��-Qk Yg_�ۣ�'z��')�Dd�E�k��4�X!����o�)�����:���5��mG�H��
{1�]
�d$����{�9��Z���X����D Xm�T{2��y��$�F�䛦�JL�t�q!�r�l��!��y߯�&y,;�I���K{#��S"ױ�S񈭻10��Fw7�\�q�P3ul+k�>g����a��ѓ*j'[rmlw�.`ت�G�1�%l��6�w�#�a�Gh,G�������[)@?+~%�����c"˷�ֈ�,�j��
�7�f��s5ﬖj?�����Y	-���k;��-`0<�K�>b���N6tP�foE�ܡ/�?-���{u@���hI��p��٣j�*�Vm��S[b�4�i�����Qe��A�7��(P'y/g X���Y'D7���R��}�Q!"��I�;�����fZ��$�	9���d���NH2�&V9�˅2���V����m#�
��;��GKߛ��1�7	�}y4��J-1���K�x���?���_=��^�3�ƭ�K�K?z��!��I�F���ѕ�4�o<�:��^��4Xщ��b�W��ӄ_f�v@j��9�G�@�����l�ߺ�	������ߴ5�Ba�e�T���f�D}��ʑ�۞g���/���y��IW�Z�&1�:􍒧2�̟ӄJ_��e�gs����{�!I�x���=��a��l)jj����C��e��o�a]c�܂�����$�����j>I+��r�^�T���'~h>7WןK�Ap�S�AA����2
���+�� `��� ��i}� 'g��6@\��8}�?Z�����W{�aj���<{-`Df^:��ߗ��GI��	�q����OwcQa�%%%�G�?pk���B}����'

t�cQ��ז^म/�I�����	�X�2}��k6`i��e���l3
^Y�u���J�0j�G}��ԣe�|�轞K�Ӓ���T�[���H�kk&A>>A���'����l��m�xd��]6���D/`$]���82�Ȃ��-�_�90Q	L�,#o�1!F�		��4�r4���jjTk �B z��G�<�m�p]]~018�K#{z0�wv��b(��>*� ��3�z���D�K^�LN�u���L��%Ɠ���6���_������w��ō�������Pw�,we�M�dX%����ꞆZw�: U��c����ߍ j�6g�V
�06W8N�Ե��EQ������{�ը�z��6�._B�l����<) ��-��VV��$w��y�<=�xEY��"/wq����?�ћ���S].L�s���E�ҳLt�m�s��]���cO����DH FG�L�/�`*t�+Ͼ6ӑNf9Qa�P��2v1�E�����������un|��,�{˫K�ʦ?�(���C�=w�Oeeè+p����D�Pp�O������%����ܢu���Q\��#�h����qP��H'�I)����F�F�,�[w�:�����s亞�?Q?G���:�˝����9fy�h��n��ν�n0�+ܓ�����ɃN����l�V�_��dؽ��'��G�U�wCTB}��e��6�9ń�I�E�J����;o�c�%l���Tm��y��!u�Ն��e4��ղ���|o�=iȓΕ���QQC��Y����I�o�c�>��a܈wݳ�N�:&|n/��a���#%����P�ۂ"k���x��:/�\��|����������Gs^�)땼��[u�)j�FM�h9Z��(���|�������!i�$�i���B�˙d�Ϩ�X�X�g����_T�9�^ڒO��!�Zt�v��Ǜ6��������ݧ�V/S�Z睔
G\�F��J��9�*ԏ�Z�i�fo�Ϝ:>���F;w�u�<��a��K���c�{���T�6!���e�������\U^�G�+T�
���S	��ieͧټ�aŧ\n���W�u��'�Ss���7��SP����ω|���̩b��������lP�t��-��S��7����gf��|6Hrf��a4�/�)V�9Z�!go�Ÿ�1nf���G��-=�0��p1^��A��к��`<O	w�O������r.�MÖ��0%���=���*��Wݵ���u�̘��Sՙ��Eg�EQTQI#3c��S�VQ���UA!�C�ִ��S�,�:$J	��S�cJ)I	�s��I��y�6ϟ�~���k�����}�}�{���v�W���z���������<Y�-(�-j"~��!����R����4�s׍Ĩ%��aH��t�|�i�7��7塜?��m���a֥��9�Iڎ���]9��������v���;Hj&����Z�.mg��W�_�!�/RXt�L��'�[��k�m��ͤ��S�����"f�ػ��ɲ���o~����3 �K��������x^�W;��->��X��ן���6���ȝ_�rӄ�-I3ȅH���=Ц[p���6§ݦ����r��q���>>g��[���a%��(���j�;��qX�Ґ.�׳ܘ��̳$ڠ�s��J�ݤ⥖&ޮ�[U�'��G�_���"t3��Z[�3GFY�[s�	��#�۵����G�L���^�Ll	�V�骴�ڞ�z�:&��O�n0e�5��y=���t�+z�{X�{#<��~F��l�c&ux-U\��k��N��.�}TgC�h��� G�[5�x���r ���D3bc��4B�.�>�0�b��4H(�?�I��-��臢:H/���$�f���&�1؍F��4|��.xt
6H�����՗�](�.�#����,�y�(N�]�c箾Nd��i��U-zB����&@���*�(K���2Vs��K�z�Fٽ����֝C!w�_��m`8��E��3�ؙ�ם,��#87�)�>+�4*N�~�@�g��-�KMe�r3gֈ3����T����Ń�?[��*ئ8�ʪz[�x���z���DK|�|��ı�;�����w��q3=�R�K٥�ՑRL��I��q;Oڔ�L��6���Z.6@�k��{PjH�Hj'��s��'^�L��s��j�>s�U��Z�/�X����j{�*�6S���@6���/
�L�&2f=͡�u�M�P�E�.a'������'0� @u����s���M>�k����L����H�.���TKnEQ14ec���r"�� ��8gd�y7��ykkw���0lΙ��7��~ct[8�&,�59m4��S[�Ȁc�n��K6�-3>�ٻ�|ҋgEԣ�I���������0 ]Ac�Y�и2�c�\n��@��^ ]׀jn�W�$ϓ���Z�5��e�1����)h%��d��$�������Xo4*��k��N���N4�U�7|�H��tȗ�}���|�p,ь�~���z��;|��]����+8��		8a`�L�EQH5�:
;�`���?+^.���<�R��~���x'�=��~a`>��Y	�i-O���lPE}Vw{eV0;�j48�f��A0�l���l�k���?O?0�؝Ѳx�|�{��\��ނ�<ؙ����?���4�q��a����V�Z
���a���N$�%��Q:��~Vl�����l_8�=<�r+���U�]P�����e�c���|Fvc���v�hb������2g]��s�`�>�S�$����W�{_KcU@��fǄ����9Ƴ�jG�I��l?� �qi�X��C��Wϱ:!���V=]��7|Do�0y�|ͳ|5��HI�X8Ӱ8�=O�G����2�a�����m���������b�Hst��vIb�Ѳ�9�C��'w�'�P1�̘�R��rm�٭�<�
'DK��	>IIYY���Gh`jC	��ղVI\����H����<~Y���4��`�w�]!�t
vس�%��N=�zS�����I���e��k��hci׷�bI
���$��z�XӞ��:5̠k��G�U.UѰ�hW���۬�q3�������n���h�{��33җ�I�W)]��?���5P���)�D3�Y�a�W��@O/3K<�������s�x��j�g����6���NL��E���2�U�\��<�k Wm�q�#�>�(:�ҍ
=Shs���l8+Y3�m�ź�+͖7��NS(`�D19O3������u��Rw&���Ly�� b{َ9/R�C/ۓ��)��e����EV�^f��� y7GP�R�3�!��"��F�1�q-S�K�ǩ�����I���0`����g�e�E��ɝ_��?-FI���ŅzkD;l�f�x��D���j�!����4��`�I��L��fRX�^ї~���[x7}���-D��]�Vr컣�	mL�[Ɓq�5�V\��j�/z��#�⸁6��O�X�RS4Kp����m�|�C�5��/W֏�����fZ��v߼f��OVG�>�"�5�i`��ͷ�`s��8P�)>���VS]�*����|�y�94��Hz��w�ݐ���	M�ݍ�w�>9P�'�22�g_Z��||�	(?4n����1�A=��M��{���b_�����cBӳ�h�N�폯g?�+%��Y��G)�D��xC/�PA�e�C���	���`C<��H[K)(��H�OٜX�S{�S��~1�FW=�IƯR�E�lg JZ�0��% �+i�koL���G�</Q�0zy��5Ѵ_�b�9jf�5ð�L�o�n~�o��c�߰��z"rs]��3,�mZ:7�������Fq�M����#J�gg8k���={-e��0�C�f�Q�[�'�$_��\>H�v{��0������\���!����S��\��*��Z�S�?@:�jm�L�0 U��ȯ�{��P�t�V-�T1ڟ���Zp�l�W�(b�&Wc�����0.g��Z���dӼñ�ѽ���ʮ�F��;�=��r�T��P��Ǚ���
c1x@a��$I�+3AϏq�ځo�z��Oy�\�:��@�ژ���
 0����mG�1���"S7����x�],єA �W��3�f�a�xA�j�0yB��k�^������2�V�x�	]�����
��`�+�� _��E8��&�΄��-\��+������S$�l��d�t#�
F]�^�k��	!�X[�V&�[�PwJ�vCc��D�o5r������]P~��cd��\Ei�}��.�G�
�D�c�~A�gD�����^�X�r��~N�k0�M�KH��o��"1��iIĥ8�P��P��'\���z���Y����/�A?_�*�6jg�l����Z~���>J��0��҄{�����A��r�E
��������;u�kR�b��c�r}�8债"h3��|�դ�r��⢦�z�:����PU�6_t4q�sҫ����!LSt��+��#�Z���� �������_�;U���!T}�ϸ�2�,�R!?�0���M��<w���³T瀋�.���Ҭ�QC�6g����|��h�F�gSs3P��G��e��e���AD��e�х��%XV�tq��̑�n]���o:._�tw�X鍛ԏ��9���I_��-��#�}�Fk4��F2����m���N�p�����F�\��_���3�;�vF<$�8z�*��K�$�����?`l�\�`R�nn�t�zY�4��aN@��B�r㬵�j5ƪ,�Z�_+�a��{�s�N='�c�gE��F�mKH�sٴL�6��.�rO�pO[�D.�J����-+t]�K�χ�k[ny[�
�߷}#�+RX�C@[�Q��+%�Рy&�
2�8d��и0ʢ���k���Ȁ���k�g��=������������ D����_jIC�all,g�����t8�.M�&+j����1G�8�������- 3j���@�/;7�=s�)~N�6-�5!�)h�e�2*t��%��!pZ٬
�����/�ggo��=�x��/�k��X̴�zܐ�>���m{N�K0�RI�IaN<Q�GxB�W��r�W]sK	�3��G�#�.����oA���G�$�:-x�v�o 9��Te��rb��R�n�
�d��aQZ�ܬ�(�1�/s갼S'hޏ�.T=�g+��8���"?P�r�2$�C�[Oŭe!a�X5&���>c�ﯟ�+�/�p�;��,�?:H�$yN��a�/��T�]:�>�,���\·�'�ͩ>N��?��#c��W.�*Av-�"Zw��r-f�J+�|$���+�0Ƴ����g����� 
#��/�/���.��E���G�i��A���.8;7*ܕ�6|�[J�-:��7����y0{͒�@ >K�/7b�uC�c�d✪�w�6o��L�m�/ �~�K:��.4'i�}.���Ѻt�Vn�S5ΉY��QZ�؟��+��eT���K�+����$7���l������L��I\[@i��. �ʝ��DX�E����p�}��|;k�E͢�G��h[I�\
329��n
���BQ�u7����Y� p�t�@7cz�3Z곱���/߹ �HC�e�������g��w�y���a+ECqDckݜȈ#w8k��hv!gS��t,�v�Um 0x��i&�zt��?.��g�f��%Z�f8�� �s0���Si�3�k⁮��6�$����LQBr���+_�H�[22��6��Ƿ�YǀмЮP���ۉ/�J���7j�{�����T����_����tns��I ����Ι���P
������?�>s��Ü�H�@`m{��V��y�.�q����ݵ�OՃ؏ak��
���G.�o�>��3.jڶ�R�i���R��3'�(�q��?����06��ܭw���_w�@Z�(�Ơ�J�5�-[N��]���9����R+���Y�ݠ�q&w ��׭�q���_�🞣oӈz~��͏�!�]���2�X���n+M�VZ�O+f����m�-']��:&Dq�>�����Gf��L��N%�O�G��< �g[ ��h����) #�����E.�Pu+�*���3<|�Ku)i�����m��Q��Zv6;��{�	��o����֝@�w�F��cu�
�d6?1���WX��]��PM�M�L]�j>S�v%�(D���3v4�s�`� �Yկ ���99Buf�E��i���i���]�h
 ��i)�"Q<]�R����7�|�M�Y�;���C
�Am���zDB�1[��#���z匚�gs�������b@D��BC(K䑍��h�~~�н̝!+ ��[�fĀl����(��#[>���lq�<V��-< ��-Gq+�*&���a�Wmw���P;2?��-��� 7��e�Xg��/6ט	O
m>�����;����X��@ �y����[ ��v�^iJ�kPh�����U]<��K�08V�tm~,m+~I��f������Y:.���R����P�����f��h�WQ�S[��+ Ͷ+$8�v�S��l���%��V�%���ԝ�1!l�m�d3���ȇ�2F9嫶ߦ�5>S�y9?Il�O�%�KX�C�w�3����4x]�V D|����e�Ur���~sN�CBl�ɼt����Ʋ��t��^��B�Xƶ�)�z��K ��� ����Q/�+��S4�w��R[�����b'��,�5mb����W�^��p�A�C�eU�S^0�w�Y���;2e������\��2�6x�_����#�QY����v�����x�`Qq�.�̕��55J�=@�{{���B��'��'ߦ9��I�+ilO�I�'S%?� ��7�S>V�zU ��*��Ƌ�wt��u��$�$��g���J��}}�]�G\���Ñ���O�~Z^�"繨o��;�;C���I�2�+��@�R�8n`�N��Mſ��Ys|�2��t'��5W�M7.^�w�G��Y�eD�A��K��f�>{'�e�8�������g��ϡG~�����\�N/��	��{���v�-r���`a�y�����$k���e��z<�&������;�K;�rv�2��z��=�
�$����7�j
�C��*_�y�>�\�ӆ��$���疕z=�j���}�^ȉ�����3^�\������t^V!>�S/��0m�/�����e��LX� 03pd/]~���(���Pv�ɮ.�����|�9��S��j���]�(�J�{+ES�߀6��i4u�zw�+��^�"j�� ������:����[�:祦�E�z�6�����u���m�]�
 �y�,��Q��=�Ӗ�����R���EL��e�?l�#��{�PK   �v�Xv��� f~ /   images/4d249bba-3190-4770-b321-fb8fc027a237.pngl�	XS��=��-��P��(We�@�U���2)a�)2�\�N�'"��@9P0̓��0V� �� B � ��oZ�����<}�޳�~ǵֻω׎�Yl�z��[1��9HH�TKHl	�,�䧙�g�|�+��f�O�f�����ly:TBB�9�練�'�*�9��F8�-A t��C=�{���f��A�ۡ����辱Â����{N���N������-Ү�7�g���װ��6���������7!AAQ�}�C�����w4����K_��������R�{�����j1���}{k�<��=1�VF^x�/8o��P�p�[L,��^Fi���0UX�����W�C�ʰ�e9�N��'�"�1����J3�����B���Y���@�ڌ6Fն|/e���YMFb���7Q��yp2&�(�0�6��j����Հ���_ڟF�Ǡ�����c�t��ZD<$����}��p=�bu�l1|�m�)L�N�Z�ش=�Qm_}* �5�)�6�dK�.�
�}s[\�g���L�
Gwj��Yb�>�T�n"X����m�Er�$	F6��fw�oV�`r�������AU��b9��X��E;Y�{��x�nް�m��C�qF��p�8ƽWW��^�tO{���1����?
�1�*b�~��wң�(VN�[���i{������ ��91��\�-~�sA8�O
���R�x��BL�ġGgº���j�� <��qx�V�{沴1��tfo��qҀ�aHW��@p��H��׳����*x�
&Έ��X2����]��;_�O6���P�Z��D_;j�g�9f�몫�fQ�̩��22s��ܾ`_�?���0H;�Y�\�ЮB� W�?G<�-
�ѫ�С'�$K�<�lɠ'�����D^��@�P>�p��9۸�妡��(�n�O^hb�^�a��:�*��GA�0~���A�̨��r/����
� ��T���R�>�z�
��2��7G�jL(�PL-y���J�#ݖ0|6\�ѝɒL
��/�=����FZT�GA�`���[�8-���P����B(���0��+:���%��<XǞ��F��ʤ֜�����t+�&<у�R��(l8r�9��~�[���@r��2�4Qs[������^J�+��s�
P�L�|�H�$t����Gl�5wZ���v�]7�௠�2����'��|n��K�NcB�������œ�=�O��7x��̹v	]�+��6�ryS���i(f�=a!Yx��b�;�퀖3Qk:�����m
c��AV��/gG�,��WQ�e��^
(��WupA,��}F�o��5�()�75�t��r�U�eo<I<�s7/��a؍;:�-�J��c&��>��:� �H�ys��q�5�oO��Q�E�1�h��h��~���p���/Lg48'�����yb��J���;�70�����Є�8�)��G"w�\���*��á�|<�1��Oq���5N�7��3N�	M�	�x��wJA�I�AS�_{�ǰX�4f"&-�nӒ��Wh7q�>�\,�z?�Ҍ���:�
���M({,\���-��\���ip������R+np�4ބ��������
��(�Tj	O�D��0���.FAÖ!X| ��(|�cA/x¸�bt(7��$v�'@���d� IܑUYZ�<E�F׬|�5~_�j��l�$��p��l L2�$��M���U�#܇�Z l;O�aV�\�e�p��8v�*.�-ʜO�%�t	��bA�3M��s7A=�	*e�&*�d��c��P�s�4��w � ZJ���2p�$v��ʵ/�'��QP�N���y�r�S�$��6�(�{��)�Ѣ|�1 ��"ju�౓؆�)��q��	��!�fd<>�B,�#5{�'��}S�;��d���B�x��~*���۲4�*��%�ݟ��0puEb-�����}����,!Ḡ���3jA�X@�{��9ǰkA��_u���C���Uv������8����^b��`���Z[{{NFN�����fR��M��A"
<p��O�̬Q���@7g�C����L*/���g�Ν;o���<�x���ӧޣ������fM�7�.w��$��x�p�G���e�\i�T��=��-��L����Km��*���'��m��t��Nc-�O���0V"���&����������Wd�nl����j/�~�����Y 02�s��]*����E?�'CY:ї�)�//'�������K*舃��mɮu3팆�t9��\R1Qy�nv󐁢�*p{�>���=J:��a�o�S�ʽ(���#0.� �-�����F��赶�֯i\L��h6���Nt*�*#3��H��ȵ���>F]PLla��a���㞞}u�#M��ȸ������ᄞ�R5^���[<���ZҴ�Uߕ{wt��dge��v;��� �ȋ�/5�LO���I���ynO@{?�.�,�A~6u0G|�a��P�=q��P9h
ix�~��|/uf�Jls����p�%���XGz�ٯ�8��Og��C�ePG�*ãQ/8��z���0�C��>��7��6Ӏ�97>��&���%�j(q�A`L��<	k��L1]`�����}=�R g}yᖸ��J�=��� i�A�탢��^#{ל�-h@��)7�2�K��W�^e�K�ڔC;�@Q��	ۤ��1����+�NJ�ݎ�yL\>Azس�Z5��k��@z�H� d�,.x=���Q^iS!�F���ȕ����4Ǌ��:xB8�Y��&�&��Zԍ�۲I-)櫋�����<6��
�6�i��W܍��yF��/�N�^TF������=�i��t��|`F�$˟Z�Sf@��t�XY>	*n(lچ�Z*,��C�k`�=�E"L��{6[����S��
B[�~e�*�w���`O�6=�8t�!Sq�����^}������fO��"�I���ΈuHޟͱ�Ep�mS:�#��d�F}|h
��V��o�/�SOF����8���$>���Q���l��N��3#f)'��rCe�9�Q-��s馧`���)&ô㜾�tHE37����wS[�&*�cJm�x�MY��}�cl��7�E�����b�A"]�.��^!��f��d�d�����Qը�2nz{e���-��w�`�s$z�%���E>�qP�w��y����d����`V^�Y�D���œ����˙i����| 7�yy�"h�H0��_
���숙����r�C. X�誀3��$�6Ͼ����R�i�ho�c��m��ZsKQj��I�4T\�$Pv�ހJ�C�r�jζ%��7p�C�<���.�㥧H���f ��AT"��`~�ސ�O�,��Pw����[��6��ͣ�
��(GnW9b�����T_���}�=�������b�� ���ct��2jؒ�����U�cDW�pC����$���c�A�[���ױh7���ⁿ���|k��4�&܄�@y�,��s�*w~�_(+�X�1x��$	~��=�u��aXL���F��;��j��&�I;�oj��ωf�D����\�3U#h��S�s7ܗ?���Eb���(5DaIf;��}opn<D~����D��F�`���s��s.�*M�ܺ�BG_�
aۺBx*nP��ǰ�4kv!z��u@,�(k� 9�/���)�#_�..m����2;w�;�L�uT�?�VL%�<O� �jv�"�J���r�kS��-��X,��a��s��%���s�Gnl�f�]�,�K	R���#� Y��bV#8������ќM�"�L�C)�YX��c��lT[�/(~0�L-�4�96�VP��-Ud�7Rf�9d`��߽@	��+z�_?:�;Mq�� f5DO��$�=b�v��ſ�P��KVA7F�����~��T���2N��~�0PE�F�O�췢6L����<�nw�Vr�S�&W�ϑ���^Pa�Ą�sR�������jf���j�<�p��(�'�4�Q��zZ�c�̿X��F��7[q�U�~@t����w����$r���=�S�=`�. �2���i;W�7N�wD]q�����Tz0
����O�0S6U�KQ��j�KjQ �LP�17�|p#��L�ɏ�@=�����?Pѹ^�� ��b�޻/8�0<uS:E�;Nw%�.�u ��椝�w��3���MI�X��h�L��t�)���i1s]m����F �C��oq�F�9�qh}J&�s`�-P�N��Yw��'��YOM��y�/F��� ?n�KŨ��=[����*-�?M3�+^Jb��$�i�����M��u;��~xJ�`'�o����������a�3���2��R?���������#6'1�"<|�:�%F�`���	�h	Z;VmxC���#rbR��O���4O�3@́֜f)�?O�vm%��Ew�#�����ϑlQ��9�J�&^n�_~����G��$�%���R�N=����H�6.M�Vt�������|������}�#�4%������XC���@���P�뢒�AMӏ�2��<݋sv�⡬�:�f���%߬�� ��*��b�r�N8���7/{��I�8W��r"�3�xܱ���ίw.wH�|��G�m:f�LH1���F�.��]�3�0:�!>ÏZ�ʽ��J*�~8�=�ο�rB�G�}�1��%��uci�v$z���|���ypq$q-t��V�O�րB�v�9���Y�:��>�VyJ�W173[�ĆG�g��YԺ��S�a�
=f�ik�M^��'�\f,�ԟd�Z��	5=ͱ/I���b��8�|:�.(���(��v�E����\��XҶ��ҝA���Q�d�j�D�:2�x�Ǉ/�ƻ���e@�L\�t'�=R��eN?��LX��͉l_f��_��]+δ\��W�Ye�Y�C�-(,4��7-�2u��5Fż��}�%w	e~���# Nt��6.�������NS��wM��:4=K�z�2C�5�Q�_�4��>hl��\\�M� |�2�����U���㙺 	��3�qC����j+Wz��W��F�B�@k�qCC��|��?zX��y�_<l��8X+X���u;���!	��|/�~�ƶmۈ��[C�����)[�ϊ�z���̹��8���KՊ�@5��Q[^8
�\baVH���XQ�a`X��PE�����t��ZrD߇W7̣�ˁ����&2� ��������sZ��.���v����TaHQӈ���,��$�J �zМ�P �ߢ�[�}o�io߾dh������y�����ϰk����N=��a�29J���*�ts l8�(���q����!0;��E�ʁ�ؙʡ����	�I����b���â�~���/E����ViY~
ls��r+�q�ن��  AT��u�"g{m�&�L�?C���H�{��6���j��:���FtB�ٙ��D�|#�fw )�Qmz��8��afp�0&�Gʫ�h�	��ʋ��)�JY��Ճ�΋����[���k���i�����֤�*Fk@�gmA��{0?
�z�� y���K׈���0Ú��68�v���61�C�c~��c*�'�n��y�FK�ݼu+�2��e(��u��3F�nTcO{(P�{��G7gh_��Ϟ�p�O�8z�Dό�	홹]�q��b+#�aڻ�(���k�_
���R*��.���G��~�〴�(��܈����^G(S�n��M%�젩i��˗/��}O���-t_�vm�SO1�>3�عx�"�?�o�4t���u�D�Ak9�KpT46���,�UY��[dj�����kY�mО���TS:s� �Z?9��oP�1r�5���;�ewLw	<l�� ��6�(�x��L�����$aإp�So^N��5Pw��7�Q�������:bL?���D���vgݻw�����o������)� �5#�/�F��|,͍��2
�~�c��d�;�/�w��0E>'Y*͡�i�d��? �k�N�
'���+dj�9�ɽ§��w��a:�@X�j�+U׵��z�
Lz|Y�B^�'4l�eS��M9�l @�@��וz���^l����>�Q��o��B�`w�b���b��2�[2zf���^�L&�\�{����[��d�����aܳ��/��>���쵈�5�S���d_�:�鄧��;:Db�^K���])C� �~_;\���k~
��X��BOZ)���ĜB�6��whWMۖs73�|�Z[�^ ��lfH�L���;��H���tJ�gV~��dV<���~��0�%>�WL���kV��FIw���FO�+�\4��M�{gMF#��cfӑ�S�2���7�^ݺ�@�����"2�Q�'��ǆ[q~�}Ip.�'!��\�<�n
�W(9]1n����&�z#��PB��y_� w����Y�^\S{��}��B��u���=	�̜�{e�cP?��z�k]��B��g3���2�5I��L�\�w
��I�m��|b�Se�Sm�~���O.lB&4ۼ3�sW��B)؂~y}�^�S&�b�΂�RW�;��|�ra]��i��r�k@�OQ`���"�;�I��&�4H���ʔ�_?�]{�L�1gϞ=S��i�����5�)�E��c&��dcgɵư���84J��N���f���Z�+A!��n�|˼#��n��O�<��}TS���YY1�g�.�V� 1� ���N}��D��5J:8�;� F�b,�-**JW}�N�OjQ�]�p#���x3���j$�A�ry��L�������ٗ%�- �f����F�c?+���M���n��:�U�L�	�B,��fJ	Uڌ\/	2����u��bX<�^<��8$�I�:��n�n<n��%֏C�:a��	�O}��%��G.{4zrL����C(��>_x�+��\�%��I���;n|�{\���~v '�Pz��{��޺�۸؊3=����8w�.'XrQ��p&<Յ%W�o/�c<G̢�_5ǂG���+�yV<��C'��[�f��{������h����*U���o�F��`���ͼ򷙼D,V�ň��d9���^�B
͝ȼ&�_�w��	�\/�F,�	�g-�0��}�di #��>�WRW�3��irdw�H��#+�H��/��N܀��R ��b��(�VG�V	I�y�z�{l��K�G�5d�ʟ�_�3��Y����Co�c�zz��o��Qڈ1$x��u#�C�>����t�4�5_�������526!�=HƯY@k�6����';��)�b�,L�il�VwZE��[O�3��g�7v=}�tkϧI
�<n����~G���΀/@[���d��1�ӈ�|�.S�9bs�`qp��O��Z?H��\/���I+ŀ��>��FI�3� ���`���1ڒ�z���`�.ؠR�UC�й��.�+�@�'����	�>��.v#ԸSV�<�q� ���S����uz��X�{��v]O��f�Z���=����%���*��Щ������������e���}��X�O���f \��+U�:WNw�������в��v7�im1��r�CAq���d�ۘ<ώ<{2Ԩ!�w�ͅe��f��ؤ��/�d�K,y��9u�=��hl��G�t�W��|��fϝ��`�k�`�0��A�l=�+v�}�6����'�JmJ��+U��I�q5	r��E΋�z4�*\[w�'}'��m�o��U;.���:i��$����{��'��w@%��q�{1�s�oL,�Q��s~#�s=�� ����}et�Z�Zw��J�?eKa�2���pGlC�}!Y��$��t!�G���a	�))�������\��~~S�7SRxv��wPj��]�V�{/��`�-�o]����H䅶�]	���DZ�f�;E�h�����:>�&����8: �I�c�%��0��0:%C�7��c��Ka�Z�0qY�/y�8b5Q���j~��Z�h'��!7�%��M,�2�簈��������S�]�ČRC"�6NHt�:�Gzr��y���rA���
�C�A�ȈD���,4u�����e��w[�Cw�م	,��}�b�����`rr2S:�����@�;Wp��#r�l��O3Ж�cF��ݔ�x �����֔V�0/cv
뉬[�=K�ӟ��rҨ)�nXM1]kt�燌Mٱ�P|/������j8p��&茺�D�w���6�(�4�9 �f�#�k5��.
���^����j͈8�f�����B��K�̓�=�v�\z�R+���I���v�7��a��-$�^S�b�*}����>�&�E׳2��%�62ed3�0�i�51��i�Ob]�c}?�<���䥘�>���}f�	�}^n�B�n��o@'H��Dq.�������`x^T��@�?���yϦ�E�vj��q/�܋W��Bb=� ��FǞ;�r/��gg
�'��.~I����k?P��LdVN�eB��`��6�R���K�mb�f.	�h_p<ΜȌ�I�p�eJbZ��$���Pkf�0P�K�"�l��n>xY����^��Vi��l���6.f|��Uf�]遗���n����/��͋���0���r���Ϋ�1,�d��{�5�����+��[H�����		)'��/��a����r+C����ġv�"�������}�0���-�)�lKfhU�� ���r�j����	�]�W#!CD��a��ń�l��D*�J�=T������=&P������U��ow��H!�)O��Q�Xm���|o��� $VQ��ޠ��b�Z����/:u�C�!���[�4��^��	��:�mE���7�H=��/���E}3�J.3���;�Y"�^�R(��7����zP����j9G�&'�r�
.5�~��
�������{ٲ1�L'��[ųQ�V0��a�(�0썝�F�ڇ8pT=�/zC�"7�N[���Q��755]���
��{�]�F�ͻbK��۱�0�
���NK%�����IO}mo$��.���R�k���|��LO�����5l�0Z*
����wPN���%n�����g�=e�tP�;�οv��mz�j>�a��bx���W��®�@h��o�&�۱k��SX0��b0Ă�L������������e�5>�7m���d�ơ���>�34Z�Ʉ�r�fҿ��f!&|�Գ�~NNNW �N���0r���<l_����'���b���!Z"�����b#@l6C�OF\�*	�#�c��P���٣��p��K�M�a����]���]�1&6�X��)�-�v�X�6��r��g�]���Q�|:v�>c�'�}5���(w[��-CB�@"�̖[� J��D��j�%�6�kn���a<�/v~�r�ޚ����U8ه� 2I�.Ҿ}�����m �9�b�D<�:/k��/�EwL�!P�|+���A�sJ`)�� �te��);t�frՔ{���xjZ���shttt8�r��xr�v\g����<^�ܰAv�> ��n���7� ��o
��H��mL�ڶ��N�30�����aml�3���u�]��(H���&ƀfkx#���.�Ef����i �Bw�@�?R& �;6�V�<�����%x�����<�M�L���1��w��;�JXn�uA���g���K��Oa;�,��~%��#V͆k	�h��}�\�c:�j`XgJ��D��_�tu����%ڋ+2��ȉ���*�Z@>��Ø��2�h-���1�g 5��_'�jFt����̣	j�<�w�չ��T[�_>����:`��w�~�u����@⯵�;B���FW�8dn����1U���R�/��En���
m*�w]�r���հOnq���?r
����x]���Sߝ���yݬ�nS}j�r\�J�͙��;�C�Y��e$��!��8�$O yݼ	L�F�;����x�ꗒ��z���~��*������+7{x��s�0�?�+���b�<ɭ���2�=T`�F���C?YB��5�¡=�V���Z3���E��׈���&��҇]�j��z���0��R�
YulX�J��!0�H�z��i�O�g������{*m�ּ�M@˟���bʟ|�W�cV`.V|1gOݒ�%�(����3�B�7�U$�C��w����5�Pi�u��
��B;�5i����M�L]ҙ���������������u�@�s���ߤ�@1f�y�����5~�:�'}�탕��F2�KS2?5�$�oO����9C1e���̎�L�����f���O�;��g>3��jD���*:$HQ�yp�;	�IK���5VJ� ��{[��r��_P��d�͘�:���'��d___�4����19(�C�Ńhʩ	�^P1�>/��P���;$y?����1��yq=QԊ�[��=;�lb]��������N��%(��LA�E��Q�J�c�}�i�\+�3��Ä�z��
G�����au�O͒Rl��q[x9�6u��ӽܡ2�Y��]��OR��-]B�5�\��X��7jrU�8<2�hz�BGqv�+Є�{�k�z�\�2��5�ĲC��Y�:g3Me��v��2�,���Ĺ����Kw����H�var�x�!_�7־�Q;^ߏ�-z=�k�L���D�**U�����VZe��<z}d���xzK������cv���MgY���d���\�J�}|N�����~��}w�cφB0co1�	�Y����2cv�Y���K�M��tp������j���I*�n�!!!�D��kmGH�%<�E5�f*���m@���:l��zs{�y����K��0�ѷ	Ԃ�('�'|�+)<����g��Oz��5��e�j嵅�k�2U��� �_Ǳ*v
����^#f��H����hN��PC�#ƍȤ�X���@��vIp�$��u��ܧy]9		�"s�ZO,&7�RM&B��<w�OM�e�L���m��-C��4,��1��&\�k��]7$�g|T5~y���N�n�8妀�����Ж8��o~�dovv�­��㴋�K;p4���n[^F��%�:�=��H���yM�8����YZ�ڊ�˗�߲P���yyO*+%��)�Js�%��]��6_o�|����MOn��L�����t�ȁ�EQ�x��{�c���E'��'IJ����-�ٍc���5T!�=I�:�5��}�"E�밼�����~���u'�I���C8Qjvy%'�M�5�}%��|�z(�?ȫ1��p�mb��$�}D�$o���]�����Ę�q,�m*�Fŉ
���cIj9��s�j��Ir*��֛$�b���0!O�Q���G"Ӄk�6�4���<Q:�3�$`&;�I�4��7�ԥ<��#������)@��?yr;QZ^�oT�1���T�CY	9�,�"4q���Q�ר��SQ��??���*'�p��;�	b���SQ�}
�V���{�n����Z�[@�^���֋�,*:��=���/\��.�f=IM�J��{�>sÆ�qP��E^�J�[8���#���O#������D�Yq�p��~��q�6I8���ar!�SǪ�'qo�x�l&a��0d�xJ]��cy�jl,9�HA⺈dyW��r�ti`R�h7����������wČi�e�t�f�&�t@ZN��k�4�Xہ�1�H݁���X.�\u�RÚ��]�ݛ�bs�&��ƀ}�*��͏)QIޫ���i�Y
��O����V����@�&�A��9���4�c]d	߈M�$8���fh´D�-�5n��hK"�d0����>\O��m��Xl툺,�2]I�/�7���IB�%B=�z �$�p��0R�NI�+Կ��bh�i�ǇIR�h	���Ƚ�L5�ɫ"��Z��|^kf(�l���	������8��.ryq�/2��?���p�&�w�9� �R��`����.��*{��Y5�/XM�_��C�*��$����$�覠���  x���#f?YiI�Tkex��;�,�b����zJ�)�>�M��I�=�^c�C�hb#�ʂm"-1"k���G��ʊȫ��q��'~u.����ƍ7����]A�զ !$>�J�l����0�t��O�����~���Y��r�@>���Rjm����G�~mmm]-	o1l��E���."W���8c�MC�p�ed�w�o&6i�$O���o8<�m�!V�m��w���Ν��/$�?	NB�Zci�.ߣ�Y�r��J)QH�8Uň�#�A�5��|�z( %=�����r��N\mxKU,�y�=���v8I���V��R�'Rq�x��|�؈kp���4N׎�m��}#"�S%%<0���߲��Q������8��\!����h�V��m�6�#ݦI!~WK�WD���Mݴ��*��ȳHOs�$ʛ�3(���d�K�?L���Y����H؏�d%kV���>Í��>���|��7�I�B��űv���B6~��|[��q`&�*��6ܼu���\�	�9���<K)!�=�gy�v�&{�3g~D�撤t�q�7 ��G���~�&��NR� �%��.�b�A�&��ִ�m��`���C�Y&��:Aʈh���n{3`a fՖ���4rn����'&�>�i�"dnǥ:�;��v�Kޝ�'O>1P������{i�S����d��[�閍9���������̝�+T_Ϩ(װ�&*=-��=4"�!�T�2�:�T��$�aN�����٢G`#����<$��L�.��G�lB��-�]�T���*	��[;��!��W
��2:�pO��HC��!��p|�K�7NVEJi�����u�W��B?��FZ�D��L/���Px&D"Eo)vq3j@,7RU&�>�ΫKsa�yi��m���2?�a�Y�۞n�/�ޡ���f�ǩS�΄=w''']�^�;h!)��h�MF���_<~xc�u��ŻFQ�?~�tɑ�4�\Z�s�j8�.i��(�]��b�j1��*�Ӗ�-�b˦�>˛�Ns(�$��˽;�?C�5�R����Pd�(�겟�͗?�������o�$Y3׍���~g""=S�*�y@]z�c���Iv'X�onnn�Zk����dz��545�%$~��h��!�t��w&�<��u�Z�C����r�����]i��8��� �|���U���O�v,	)ֵ�]Mv����W�\A����ݮ��<�U5 �!�N�c�Iᶢ2��'��	�c�y,��wi��oh�N��#H��Y�� ��V�oDF����V���Z�y�Yic�����V9��D�ѣ��
v?���;�x}^���J>��6�|	���QU"���Y��?ۡ�Q��S���\���G�m? s*=��d)�;�w"��ݢ�Dcp�Ν�tL�3����T���#v����D�0���0o�-� G�����'~�V���x�('2[�qFF��pcC8p<+YW�e�];�|z�����b�赞�

��؁99&؄�܀���/���bAK̐5���[5��e2H�R�Ϟ�)44t�ə�>��k�= kk-ށ@�aR�e�h;v��g۪�o>|�P+�;X!����	�u-H�濔L+�*QhN}� �OL�c���X�ہ�T��{'�!��
Ę�a�0�#.��sU��:����2D"q2�.#+������*]�o��/B+#�dx<��g��OU��xO=�YN͌�E����	��

A���5�F��S�Q��������,*�����ۀD�>G��L�Sw�J?'yL��|\\\ijH,�A�&���"�~���v=�
��X^��b���O�\2���*��@���8JLL9#?J-ph��՘y	m���[մ�ZS��e����L YH|��cPx�!;Ā5��`̈́����>Fm~���\F��G7�� .j� ֓S��$!��� �����}��6�_5�EOe�`�pV��,�ʖ���i֘ �i�JI�9::�/*���֭���6�DG���w�h�� g�u�	Y��x���Ԑ�B~b�XzN|ej�Jr��{[GL��cW؋$5��cv�i��zN(LnI�sL��@��hP� d�WC�|���@�)��PU�[tOxS��,//�h��օ[�� 㝀,�_�u���.�c^�^π���J, �\�����+=}}��PUU7@����{�V�W�
��lSz��|�x��U7H��Ջ#����tedd�#h��(���Pl(���b ������R.�Ҩ �gQ:J@~�
�q���5+��R�zzּ��`T�?��Qw6�(�?=Kw�LN�`@�(۫I����Y�D�l�����BUj�/B@b#����u��s���UTz�.���S���T��>��}ܭ�����R�n`���Χ;�{�]|_J��8P��NV��������s�� ?��th7[�֜}��*P��?S����'�o�����ۋ����Q̪%�Z�J���d��'���0��֣��¨�{�|�pVN��= 3���p%p�,��?�G�c��~���y����������{  ��������Hi����b��X�@E�p�r�wՁ4O����������A����>y�ys|ǡ�WQX����� �Z�bd JK��B����kV��o�w�n�\���u-{��˸k%Ф::bڲ����_=G�����B3w_��+@�;#nݺ�`������y~��[���C�r�a��$�`���~mo5����C�� rZoo�9K����c��z�:r?77�Nk,�6X������W�Ԕ��G����$om��+A��y	�q�8�E ��a[.c��}�!�>H����D0�u��볏�vQ�0��ͯ���h�g�B�Ɠ�0�����v� ��SK�L�Y�G#�w���#diJ_��2��� P�`=V���Z7��E�oL�*!5A�s��X�/\k�G,i�K�R������	D�i4��Pz^eô,UI�U����@(E��a��)�[)���O� a�`-�B�>�-�T�B~R4��"y9	�f�)���i�	�O-9��W_9A��k-MM��8�Є���%�P�2 �ҽ�u�z��o3��VA9��1U [O]��f��E��ٛ�@��F4G;� U�yz����DϐG=�p��s�As�u�Z��*y@�21q�4�,���~>[:,A�jڥ����7/Zo�읉�73c�����k����E {r�$�h�VCړ��I�U�V�vj�kf`U�F�	�x��ъT�c�lA�1�n�3�o߾�I\Ɲ|?	`rz�8绮X�,��h"V�Ov�Ծ�-� �a���e�agg��Pe�֫t���u��9?�$���}�NG���Y@7
8��~��d���u=O�w������Oh��)v��I�?@�;W={13VG/q�*E����W('M>ɡ=@������g���u�"��;�5ѝ=P�����70f�����Ѫ���)�j�Wfǭ��/��I��-j-2Lu�L0��]�* ���	ľ�Ӄ�݀%ש�m�%(hh�*+��H7��k�ĭ�1�4/[V�!纈 ���6vv���X�?�a�Q��n�$�l@�t�իW)�5�;���n�-�!cO�� ����%	M�NB��z��m)��R��C�.���!��D��{)A�g£J� k?�������])�)���Ǖl�g��
���ů�aD�
2U��i���6�b��߮��҈�H�]�R��8Vڡ̬,���.0���7T�t���N҉��Df�H�����r����B�'�����';>������ۈ���xfcqq4�I���,P陃Ue�P`��%�cJP۵�%!R�O�4��H��ȀsF�t�Ò$k����K��~?��\�w���\%;:�C��}����2T�3��*v񈼭h9?�v8�k���sp}���~�uua;6zz�$h����M�%�{$N�DO��R�Lq��Z�v���i6S?B�lY{~��ǜ�ˏ]�x���WS��!�?��c ���G�0�1G�S_���p]�)�8V��O@�lml�� �\/�u(�~۰��o���
M���͸�Z���ΚY��YY
�������7ե����}����?���g�����|�F~*Oc�Z￀�.�,P�����EYr)VB��moVI;fm4�j��g���@��q����s_��'�˷�⦥�.0+.Z��}q ���F�(��2m�S�	���̈\ǃ���2��P�4/�;J]��A�#N5��fv��yg��?�Y+�(5��v�o>���@��m��x��-,�R�'�������{�� �DjZ۹ҫ-Ye2�dߏ�gdK����="d�x��I�u�,϶@����߲f9�_�ˡݽR��e��T��Kx"`��T��g>]����{�A�O�UkhxO�g�KOj��[f*&4M���4����NX!�QPX�<��PL)5�S�OjJ�y ��HNIq�f�#�EE� ����J�����6��r��y�왯o	U6�V�4,�z/�t@O!�P�0�PP�� ��=��F50�,�ݨm�\�%����B�	jCnQ��S;7nQ�>���|��������Pf�o����I�]��ѕi�(z��'f��i|���	�A�w�Ø��&����%b��^ ���j�ZBh��!��,��

@υ#��-�E��^�(�(CrRg��"�&�A�~���Ю���O�g�qu��m
 1l�E#o~D#)�Z&�{?�h��af�� c���r\�"� �7IVA�$+-�Ut �xy�^G���C�`�o�k���eW"�1?uP����w�T����ű�� ����|�f���*CD��]�a�/7��;�h��T@]*�;o|�o��s������#������k(}dI��`��052���c�%F�I(�ۓ�Q�k�$`�ÿdkV�6��m&$~�*dl�+wD�W�+�k�4U�������/. l><}�7�����Dy�#������)�й~��\�vє���"��h���pav���"�� ��k��^G @�`���~([3�<6����9�뮃��S9����Y��O�7B��t1U��N@��5�k�B�<(�`'  ���X�W'�]m=*��R�^�X)�f��5"��  �4��G1��ф���z��oP4��QZ��By'�Ҭr�l50�X�׀Ð����ue=q�"c�Ƃ����/�o���-WT����Iȟ?UiD�j�9�2�
J�r�@���4��������"��P�'ĮO���~��a��Q�
�1!����0���zP8h��(�a~�ڠ���=��D�O���\m���h+��.$��|��b�.v���В�SG6q���D��+��j�Y�����G���e� J�n�?�̆k^�z��)�j"�	�{�\��#U�5vQ��K�_ׯ��)��0O�Mg�Me�0�`�)7��d��{n�D�3�'aK@o�q�=*���̊Љ�0�b�!0��vG���w8D�����k�������&�^c�o:G����ˣy�90��Y���x�-�����	��=���̭��2�Z���*��[�5�/A�T�_o�=����^ ���O�G�W<sZ��o$����ǯ5U3!k�_4[��:9�(>�?ȍ攫^
��O����p�F ���fh�+��������W���^����k~��Ly$�n�\s` �@�=0��s��,�GGyG�)��mC�* �V�"�qB�Z��m���w��a1q0A�:�˨�uؖ��3�4 �/hU������ �r����8-��l�J!22^�4(Y�d+�M�^�SVHB�5*+��{UV��[F�����_�����r]]�㹟�����>���s�l⋞;\c,�ӛ}d���9��B�г�+f˃�r$�X���lV�~�����Q?YQ,�cҰ;ТQ*���R�Bv��/�yyy�'Q��0�m��O��.� �ߠ�j[�����~����1��T�*B�ё���Rav+	27���O���0�z�Y5S�}�1�L;^�3ˆ�)�B� w;���QU\�[Ā�\7��_��2����ō�T�O%� ��#��o3��ބ��ɾ���_� ��y�8�����a����DTV$E�Ë������О�I���nc������9]���F��%���9y����&��f�+�av{��������c̫�vW��t	9�E��'�~<�u�vt��x�<0D�����?�N���9�Q{)^�~��P|S���]>`$�I�ɹ�B��VQo���	���{1�/�k��3:::�/���}�����I l����j^-��`�4128�˟���`�k���@��bڹt]�O�����ׯ_�S�V5���	�CCC�	u;4QUIde��������d���zy
���p8�d�Y8El��
t��leuu3�}	���&obb"%%U\T$6]|�/**j��ډ2J����]W���~�)m�{K����p�J���Vښ��W�J�2w5���Z��Bwإ.Mܖ�i��O
��������VW�l���v�I�17][�n@F�2++��H<���N~d�]��K���c�q&>������:�iu����}��FI���eJ(��&U�k	wn�dV���x�1��n�U9%��T���c�(p/%Gd�(���	;�����wmy��e�L탛�h5��Tt^�re�⩍Ӗ7Y-��˖�l:�^���jְ�`ee%��2	�U]�y"��5{��u��J��ˑ�\���
循�*�P@J�ǥJ$b7!�?���?u>N���2<���L��sG�:�`ĺ�����E����p��)t�,e�X�H�2Z�R�T��|Te��TG����ġ��n���O��4�@a��C��P�Q�!��3�C1m�JDSS�H��*a�FZЫ��g�K�[s��4�F�RŴ勺��7�z���/�G��kH222z�4������kLyQ��(]�گ?-��KY��(���yTq���P��4o}���
�W���KPWv{�wKB9��3<�֩��|W
!q������@��}SS��
���!�f���69g�w�MHꡃ�����-,D������>ׄj6�����.�rN�y�Ǥm�>�:αa���go:a^T��A2����}�D�c
�q�����1q����C��)�Й��r%w�x�>��&�
� ykuyzE7m�@��=T��@�op����Ẩ��������9Q�}q
����l8g�t��o��$��l�����Ə�\3�&r'���ofȝ[Ӂ����𗖕���g%��,�ro�����T����'��JK�tʶ��b/�TPP`������P�p�x��d��hB��V��-;�*��uĸ���F>[�ƍ�s��z����J�?���r��>f�������7�A�nB��]����3P�������m~�
�K�ӗެ��`g�����oE�-�]���>o�\�7@Q���޹��41z���YT�Pq[|�+���w�Q˳1=Q����D���X����J\JN���W�ޮ|��,gD�?��(�ɲ��Nc�zո*dqn��X�N�h����ڧ!�Q��w����CօG??=@��S��%��>���-C�%Y��9Q�+|}L�Vm�x�8&��(la��D���q>�}��5��FȖ	��GM��}%�5����b���;����i=@��M\��Tmc#��t��ř4�^^����"U� pa���k{컬fq�&Ϋ�+=��8RL7+,�IF�{466R10�LLL4�%��(�L~���rW�4��0�+�nß��c�]��g�
��sW;,B��E�iM�}�:M��
h��}0����^�:��Ǐ�UVS{θ�T��)��w�������?J]��̉����e�D���l��ᆠ����iJJ�m�~��b�U͔��x��տ �N1^
�̲���`y�*ȡ*<���I�pZ؈���r/�����j;8���mA�ϕ���o����*���A�-�����qw��(Agno���x��VE���O����(��R1�u�gƣ���!�F�X�t���V� "�g*8ʼi�vNL'v� 5V˱����x��x7hG�x������@�eϠϹjjo_�/v���|�tj�:�����C�E1�`�^���(\7�}BJ�p�XS�������������o�/��0�2���������s555|���&f��V6pbҘ�w�v� ��@�vo	������?{�l+����E����ܐ;�'E0�y�/���{��#C�����7x�;���+�
(�H(�lg�%Х�S��u2
�d�����a�1.L)�w��j�%�U��M+q맷���WVVD�#�ܻ��|8(����A� ��N/���+R ��w�ې�n�&^��ݦϛoa~a���Ԇґtt�=<<�&&P�|����[ $ 2�^V��Q�at>�Q��N<H,�G��sssrr����/�;{�w��|��5vwo8O�h"���gA��~ӈ��^@e�`Q �/S/��UN�s��%�39 �nBn��J���;��:��)���3ww3C����8�9T͸��K��M�:�Z�ߚ��`t�]i�Hd`F-��]�cQWW7]k������x�J�����&Hy\$�=C�4����@��;T���ۑm�\P��`�kbW���7�7�4�x�.2��"	ג�=���S�����H鞞�����n��L��5�U`�a���d��m�S��o3�5��S��-#?�~�
�500��� (;�D�UM�/utv��O�� �FA��s뼽�t�ҡ�C�ng`` �Ծv�����M����Ɔ/���$)���O��]��k��nr��3��Ҋ��֒�Q��bW�p��5Y�^Y$��T�p�
y�n���;w�ܷ� �%�e��xҞl���:���E2F�w��qt����{�yB+	�ʊw[��/�?��,�0f�|E�3%�#� P�gϞ����E��1�3���|�ŉ�աx5������@�>���Z�#����u���wܤp�*ou"7�{�M��4���M�AJ��������Oʄ�л��#$��\y
-�z�����������W���վ����	��,���_
��I��ʁۥB���셬�^R��ɐ������Qo��8���1�nX�؍щ��͛�?�K�����:��W�Ǆ���nN����b6y%�5889����[�w�Đ�>zmbd4^}��Y
T�/_8ED� (N�%$$�#=}�4�r4pt,�ﴶ$�I29��n3�V%a[�E\��&���V��>Q�X�ӽ��`ue4a�;T�g���C� �_`�`�(j�Ns�Z��v$��&rbk���ٌ����' ,,-K��"'M�~+����{'����jd��ݏj�Y6�?�l���[��x"oh-���Aac��I  3��[0���C(�}�����|轠�`�S�Ay����2e�<~�]��{��FGW�RV!'�A�����!;�=�%�jW:k��8\ы�Y�񣚔@�@t�c���+�"�&b#�v9��pjh��f�o��^�w�$��������|cWX�5�Hl��9.�&���v����E�8߬+W���e��D�B�t�����!��3����}�gΏ�#��O�s��j$ߖ��o�D�-�\�	���ZX_OJM=|���w<Ӹ���o�=((�7XK��0��Jo��@�U8��P�;�#��ZD�u\�?��>�{l��Ī*^��6hN,���GM�+immMX�����7H(�HK�O������2������ �c/o����v{��������.M�Ak��5�xM����,���[�i��ɫ�iQhPVn�E�$Pr�M]�(p��p\�h��QPQ�L�6�iRS{��T�+))�a���8Y$�k,�\�ZK�g������;�*�Ht�qT��W7G���U�G��0�3E��^+P�����ؽ.d�YYT���(��w�MQ�F���*���������{���A9G�jNh(����zH���q��@�'�$�6�+��/v�" P�Zѕ��
�}�ɯ��<4�}����*��E�,ⴚv@�JJ� 
G��T�B���'�AA}3���G�s�E?i�uˊ,?pX��E:]�t8_t
�n�3�*��@Џ�͋&)l�V(���
12�"{�H]8��)�76�J��"!l��U4Bw8�y�t�#;�|PfGZ��-�z���E��"�DD6b(����A�8&�re4nn�)cV�@�Iw��H\L�pL���*�qd	H$��sS��6>�d�e"�	�)�e���!���P����8�@��
ٽh��~���P����%I����*��RQ�����E��Ӽ�Ꮤ&O���J�� �!:�Ō�t���%%�A0���l�G����ܔ��`�#,�et[����Kɓ��D������n��I$" Q��Ĩ蚛s;M{i��Y(�76��҂�C;�nP���Z��J9[�g�ys��$�&x�ʑ��E�C��gݗ�A=Z���7�)��co����8���84}���aI[�,��/�W-<V��^��n�y�51��΢���qT�/*�q�p�>e��ԕi�)4]|��&�^d}��b'V�f�-_VVW�PNM�fCk����n�)))�E�>����{���D��<y>�{J�o��8L��������Z�a��d������Y��#�[a�{�w�WƖ��^�D=��dٽ���g�pa}cjj�_]}�&֘746��Lc7N�sv����$����5�܅���W[O��R�T�KS?�+���&;on�;,=�^Yi�U��o��		��/��-�.W$�IQi��*�Rhu,U=J~�:�q�[CY�*]BSSs�c����ӭsK.�����V���7@�A=��rC2�"�C�j�А.�����c���Uv���*�!]�Ųq�iѫke�?A��[&����������θ�*�)��E�$����@���*�����Բ�΀c��u��$�i�D�Бz�jΊof���C�8��ބ&ˤ�x�Y�gXXX� �A2_���`��`�k�~����겎5dP�ۺX����w� w �Q}z3͕�&��z��2(\ˁ����o�$A�K8;;��a���N>�Q<?ڌ�F�ҿ81! `i�7���q#`+o�����.���'�Ք|�Z/ҸT���z˨H�_TTT �_�:YȈ� Y�񶎎�qqqw55}��;��:<�?��F��xd��c���a�N�-���5:hk3���}��sQkmm��\D�{�=�Up6�[������Q*0O��Yr-���KI �����g.����|�!�vzF::̀��p����Dc`�&7��z�L��@~�ZKq�� �������Z&� ������o@�K%��zO��v�D5v�(����g����ϓ��"�jI&V�k>XEM��>
��ؘ!T3-���B����o���`A��=D~-� ٙ`� ��s�� ����^�`QI���h៬�A�B2@\z}q#���At�8'��v[��I���w��J�f��,Lv3:::��0v6���x������E���6���$b��(р��ST�̈́�I����;�P]966Vܙk����P�.B+�u�Q�y�)�\���ML116.���s�x�8��6K��l%__%_�s��,iDԷ3)YY�H9w��]_?�Yo���W�Lj���)4�Q��%hC3��6.�H��b�� �M=�� �z�9As��+�m��jl��@nף�H���r38��6w,��G+��>��&5$��t���=n�_:Θ	P��F��>
�x�΋?��4解�a�"��螁ktt�[�:��X7T[>􂔨��v�JH�e�{�ZP2��V��*C�c��i�хJf�E8 J�M&����ʥ�/�} Pk�����ZZZ'��V�Gwm.h��%ݔ�i��@����P�������u��Q(�4o�#���Crj�?�4!����R�[����N�"�� �v�B�Eڊ�L��l�9(��Pȣ���\\����&0h<,!�r�l
�MT��8�7���ɀ��ז��W�ve\`W��4�{z}�z///�)��Ɖ!��h�A�"�9�epx�/�`�ʊ��Qa=@՟��}�~[�\�E�� !턷�W]N�`"tyk\h
ncf٘u��2����ũCp2��`�C$c�R�jp��8�%:��t��o	�a�]#�����.��������h���{hӾ�����xS10TU�?�Zp��Y�c��Y�r�X(f�[oq&(����x/AL+q���}��࡙��J��?,���M� LH	`r"	
R�č��5vo�v�ҙ34��08E������i�pь��_4.y���W�����1E>�*�Ϗ��OG0UVU�zqPm=MĶ����:	#4]__�мB.ٗ�l����0RH�Dq}kK� �! ��e�Ƽ-�����7tn2Q㍨�H�t!+��S(�FH��K�� a�U˷ۡ��{�dS�������a�� �����C�K({|ᆝZ�Я�$�ddd$�Ő���@�+q24>0�����|Ң�vU�����1-e*�F�{���A���&��B�8C�{Od��y�6�A�$k�ՕN� �w�����<6qS�=;�5�p�����������#�T
�ךlik�w�������#��d3���e������0b̾��@ƠG	=t�٧O���ǥq�S�	������� ��*��:r�9��kME�<8�
��	 p'(�!(nh�gv8u��~����V^��&B��^�s�NG��~�kJB���]�r����G��i�j&��;���w����L�����_r�(䏉���j�!�P텄j�¸qqK�O��6��g�F=��������넥]A0�`4��]:�t�x��IgǺA���z�����o�{�#�/pp�!$F��Y:%���V��dcamSu�� � Ը3��C"N3ҥ�����J�7G_A��U,�W�p�Ҁ�� h�t�G��j�M 2(!4V�{�=U�z%8Eꌻ����6�
k*�i���̸��ͣH�C�HZ�&g��K_b���l�TUU5]]'<����ߗg�
�����g�3e��=|SX�t.o:��32(�f��nQ=7T����		%��f�E�6���iP�}NK��yP�W���3�m��r�"h(���Ω�O������?A�CT�,?1\7@�q�	c1(W0x���cʢ���b���áw� "��٥Y��\��V�C(m� ����\�=zb��q��Q�/��ǃ�Dϳ���r�|qC�A��<�5�,�	x����?~t�E~l�GJ{�1���2��lmQ�r{��q�K
f&���@#֓];�最R<]Ũ2�oCn`H��yl�N<���E>V�V���ٞi#C�u�z��j/abbf�=Q-�0������lcG���6P0T����l]II�Ɔ��iW�	?����c��W�[A�11
:��=h~A@ݗഠ���]�yn���_���6����'̡b"x72�G8I�y��iq48]�����4:z�o���;�Z::�v��/,�]:��T�����ι��a���&m�3���J����9��.Bq�t@���|e�W�J���}"��<#>!6�;�AGb�1 *�ˑPgF��@y�:xSD�
��-yQ��`8��/#��h��lg�/o�Q`K��"�r����֮.(R�x:1�Ah 9Z���q>Q�B�m��> ]q��t�v<�������t���ߒ��M?Y����� V�����Bd�\Aq�GNJZ:�
q�!e�	Cؗ� �)(���^dm��z�s9}�yb�|��볝�vTN�w8�|�����'�R��d?�v��yL��(;�h0������
�1�r;Q�VG��V5���e�����`�F�2@6�����#uޔ��#P�28l �L&�\�v�]6GX7���:+?	�9�!>��I������QU`u�Hcvv6��{���Qȃ�Wv�3U�;��%���颭%������+�����UWG��	�6�o�����)�d/Zлv�?C�=��;bw����������X?uxS���+�|�SC�"�R��^\II	hN���{@�Q|a�؅A�I�����j�F������L=�S����}���L���1)���jW�.O�Hc|rZ�+lTz���ϲ�s���L)��V��b��:�m���2[dX=�%?�I�M���^j(�����kK7�5�9����][�1�G@��M�j��I���d�����.���Z�ۂ��:�U�:+++���$+�����7��B�=D��� j��\_T��qW�c��V��O����p��`1�b �a�I��^0�=��ȢP��[Ղ�&L�I0�5%^ǵ��7�~��%�!1An3R���`��vA	h'4�@�L��A�|PSOrC8�^��h��07���iu��`�`ܑ�LxAgҗѷ��J�`���ҁ��oϚe��"��E��%Z<z;�Su��<�0߷����9
&�m�=�S{Uh04(xW{W�-�k�U���v�CGS���E��~zn=˰w� Q�w}*��Q�������
��eTO"](X��@�`N���?��bN؞Y<��.3���٢w~t�q��7]����)�Y�h��l8_t�A��N�?[L����ڂɦ����K\�a �-���g�@�CR�[/|�1TC�3��bAae����ˊP;::�y �T��,�qu�&Y/���n�uyC�7V'c ���-^X ���ń�`�f��`3���3S�E$�X��j�c�z����e�j�۷"�T)�i���L�aN+�H���$���E��z�4�ʦ��9����mF���G��`!S�f�����Q܎��_���=di�}V"�P|��B����o1���	����`9W>�ss��1�]J
�c��dBL��x�O���t~���Ѝ�3���c�8lQ1cj~�Qzd$nL/�$DBJ����'�@oQgΞ@z����:�&��_hh[@$:�s#�v��?��/���n�-҄a���E�(y`�kQ��L\`T���6�/�:R�ܘr�����F�8n�QH�'bޭwn�A�6���7�����	��y����)�蛚r>��!<Su��uZ��@����B�JCK��ލ�����)���1aD���7�`��"�G f����Y�}�̊i��VV����`?�8^q�hw4 �Gc��}bh+=�����Ӿg��7�@9ޖ���-,("�8��-��
*?7����`s��MF��Aa�u�bkӑ�8�r3�Ss��(~ m{{A@�ʔ0�+�FX��sp��J�s]����q[b6���*�p
ӣ�%oB�N�#�>e�u�����Mq
1hԱH����3vqG�������j>���~GE֦�4���+'�	SfNNzr;������B��ނUP�����
�|!	� %������c�� Z�P�����C+Js�����"���-��in�'�m ��뾈�^�i,�7�&�B�6�މ�|��b����n�l7$f�O�	L�
4lpp0A�����^�8��	y���G�4�LD�3�)��Dm�#������C£84)ݍO�:�����_�gKF�Vzy���Z�ݽ2L���Dg�ـ$$�����S�����L9@}^,�>�}D�A
� {#��P��ܝe�%���z�IP�;%�uza.I#����,FA����[��$koF���1�K5(
4%'�����(�֢pp?�.i�o|�V$�UE�	HjR�_�p2��r`���]@�-�346��)�wuuE���䡥������XѴ_�5�ݼ~G�9x��|�|Ԓ�N��%s��|A(B��ZQP�&�]�+*
p��x��H�x�E#a ��(񥗠�A��̘A�.� ����h_ƴ=�SOwC���#Z�0��B�!��V�-��ZC"*��^�03`^x���޻��{_�sy��sg��6���PЮ�**��=F�����<$1�@x����&g�R�����D��A�:땶�w�G��X���p�&�̰�8R^3҈3�AAڶ���&=��������Tl�md ��9��NdOLL�n��7�Uc/Csä?]�x�B�-�\2?�G/ds�r���Ɣ����]��&$�/ɛ赌���������j�?4�>c�!�R
 ���b����:��ZrӁ��-�~J���U`ܝx�Yh���=_�T&�]�mA�>������$ㄟ*�UȰ���dn�"��Lp@��i��--KC�7o�D/>�&�������;�������S��cbb�^�����(��			K=O�E8�ߞ�V�*#����;�V^��GS:�K�-��-YU�]���]7�N��|{}���QVzU�#�~8~��D�2f���#�q���<Ӯ�/:���VKb�]�wN��J#O^��9�R��(u�)���8�f�j���d��1k�������&IO\��+HxC1X���|�lZ^�×U� O����YJ�V��~%!f����!s����u�?>nxv9R�wJ��<5$4�a�B�HFr�q"�㈗_��'͹�����<�#,l�ů_F��󧂌���J�_^�����mV�^�����)l7��Y��	�:%����2��#��;�Q,-��AC}}�9E���R���s�D���(:�����F����������. �X�y;;�.��E�(��� &�����9����� 8E���0+����[�>���hh4��}Tk���C�!,��9sm���T&1���<��I�}����+`��>'\�!���9���w�X��X$�e�������2oE0 &��e+(;���8G�=��P�F�al�ii�
���Y�ZM˙�9��Q�G�����Ճ�SZ?�C����w+++���#|]YYId����Pv>��R:��\"�� cmGG���̔��_500�Vp!nnn�� ����o�d6�p���b@�<���>��k-	b'"���*Vy�s����&�r�h���ݻZ��-�RS͕�냥ġ�E��K���e=-�$<����J:ndd}��r.!_\�ܐ�f$<��(uV[����<�r���b����~N�mX�	�?������/±��ۥ�����t�w�@U� V>�~R{���{��ͳy��0�R�`Y�7����[>��Z�E����r��
'�ko����,������Þ�4�,**��"L���3_��냙�<�4f��`�e萷8:�þ|�^�L{���p���p{�T�պf?�����c0��g�.������f�ıCE�o�n���T���fA�<�^��$K,�'���|^[�3�� j�`�[gfR��
D�WF����w��
���=�,y�����]���(aSuk��A�0����B��������8���5��H�����}2��q�Q�⁁���X(�R�F3�����H��066V`�J�ipSc�>�H�mu,B�������l�Ν;<�����onEɃ��x����ZJ��T����zz�.(f�j�-_e|���(�$o��ڍ(?Q�jik���K۪[I�����h&$�����`b�0��>�ty�|g��٥���7��N�WC�A���::�~85�iMi1�)�3=���X��r��X�����Ăg�I�=�{�;V<��c"���xx��3Z���Y��\�P}##�}�ϒ�k�8���LcŬPeUKh%Ði{[ٜM���X�n�3G`Q
�����_�lJ'Q�����|��.W����Y��b\F���b,��=eF&&�S��7i����V|,GXQ<�g���jJ'��gS���/�cYH���l��'���se8��
�	M��Lz"�;t*͆h�1M,.�rHH�~l'���{�?��!���ĳdگ�����x���KJ����#ƬY;f9B�4�/�7�hVh�"��?6�R���5�[���v�r�dJPv��]-��{����n�Y���Fo�f�O��E�[����
��χv�L��Q��v���6�y�7�j�R�9gBt���H����y�`��U�Mglk�>��턺Ї�7�� n]r>_��rHܢ�����j�E�;�}p��풀@\U�L���c�(7��;q��-3RlON"t�+�(2Kz+(3��sT?�߳9�B�q?��ˋ8W��i���tK❺�f�S6G��o�'�&Jy|����~RZ��1oIW��t\�}��ʧ���$�^���,$<[�l��*I(���+�1q��GM� �1�������
�Xa��={��+> @��̛��֋�x��xE�������QKX�f�5����8"3]9�)�7�5|�'���K�^����w�ry�����27�K�=ε�Z�h,3�z�K��#��ŧ�Y.5EMA�Cu�v��b�0�ЍL�ɯ]*�r#B�DU���$4��4v�x��rE]HO���Y��Ve��U˝����T�Occ�������P����d�Q�q�A�h醸Q�gƆ���#����2`-�B�����uu/�sV�a\�+�z^=%����~�\PŌ��n��%��O�J(3!������M�~`���m0���*-}v�ϝ�l�q<#�w~nn���xbe�p�imq�O��I3aAA�fK�������QQ%͗232(���C�1�HK{��ff����R��Y!�+�UB�B� �Z:b�j������}}}�P�f1�~3i@����y[;_&%-M�������sO����{���n#���
<?�A�C���&Y��h�14�F��$c�,~~���g�d�x�ӉB���^�G��ѽ���<�~�E'?�dd<����_�6�w�����3B�wI1</��-�o�$}����'�aY�����a� ��.�3"�j������!!\"�V�-3+r����dv� d�N����E:�cUmKƅ h\j����)]���А��DOu���XM>2M{�\qqq)�s���?_#gR0Q-�me�t�y>~������%�j�Qo���7�5M���O��0d��� �ߖW{-��Op�N�0��HMMͱWic?�I7��Lח}�ʘ�(wn,���7l'�	}!Ng:�q5-9�� +o��e��_~����~��Pu}[[��I3�y�t�X�(� ��|E+��e#��-H��2�q��!!3a:��`_�J������ᣚ�������ZFj211Es˝;
E�wY��ExJHT�R�Z�H|�Qgć$]=��k����3t��O��J�s/CU�c�>|+[����d�b���0R))o����y]���̓` 𡤤��I~�y�{QЛ=�b<��l7�`�끽�j��8�sxCo���;���W�����*��c?�0|?lÚ��-�ܪ�lho��;� Kl�c6��V��o��_�43��:��
���ǧ�'��K��	���{/ji��T���MN�n�z\}О�A����v���%z���=���1�%?ٝl$.����%�-�$%�ؒ�\Z�tc��=�ٌWIJK+^ĺ<�iɰ������^ ����=)�C��SU��!�#�~' "�Bt�14wt�U�=��{��=܊����E��b,_mQz���x[=�,*���'�5��5�헬S��gz�k��\��Z�O�o*��L����(�1>Cup�	�Z��su�2��*jj�Y�.��l���c^?��~�.VGS���I�s��]S:$D���1�P��{��q��o�C��c9�E�"TTU�u����$j� Ny��O�R*���c���bUkfr2���LHUQ���Y�-������X�� �ђ�6�h�,ls[9�X
uuu���.�v5]Y-p[�<ǋ#Ɛ����PQV�[��a��ߗ��i��6WW:p� !�&p��򰔙J�D��7�A`s�92�XA���ܯ� Ì�bqw��>����FNN>Z�:��s-�eb�y���WC�z�y�n&�
!ޖ��2��G|�5��F���R�&� ۗ�B��AvQ�6�h5�<z�訷8�a�A��1av���v����(��N���u��0�[�W�[��:��G\������=T��X����3g`b/@w BS�a	�G�={�bgɑ���N\�^4����qk��F9j�2vG��lI/�:�ى���3� Rd��樨�7�;�����-����n �PU����Y�9��D�7�
S���g?��1��wR�  ���|�I�,��]?G�'�{̾�O�����W�%*���s�/~�˦w�м�̃3��Z��kM��~|$l0�k�n͐����	���j�1�.]�,3S	�`=::����Kz;6!A:|��y.�ı��+�a62k��H�],&-�+�����D�6���q���>����w|��ʲM��SO��W%4f;��S&$�d�L8�����d}�`|�yv~�n��E�z���5�|+^ �g}6�:�G�
���=�sUG�4�V����qT�dFr��y`� �qxlZ��y\��RA��u�1S�6G�Ջr�����i�ή�WՂ��9��'��7_L�B֗\	����m\��􌌐�i�仯*�02*�����#W'59
�R Rï��%�pB�/��Ƹ}�0s�on�6\5�>d&R!F&��Hl�]�/鞃Zos�x�u!ܸ�o�?��x�Z��̥���ӳ�C�p�L��m�5�+�SDY�F�%�V�nt�^\�&�7��*�S����It�� ��3l����0�7�yp0u�ǏPF+�uD�R�S���6�ӻ��_�g9�](E"�� N���K�(�QW����J���<oE������
Ik���CGSf
V����P�ƶ���w������q�y�����*~���J��kkyH���\�f�f�<X���p2|ߵr�V��×��4t|����6@O��B.�`�=�'�؆A#��BTM�	vԱ�{h�|�^t���Y!#C�!@HPٷ؛���>��>���Y�Uy`ֶ����R�p�\8W �dӊ�/.�}O����1�w��u��A��ǽ(�Ӻ�~ԡLZ���`w�~�|�7�G�$P��pݙ.\��v�Ú���� z�6@���?;��-��(�� ��*?���Y��l�8]p[H���P^^~�مG�� R�����'����Qt:==J���@�wɨ�؊��賎?hʁ�>�wH��7��ihQ��`��U b���7N��I.��
�
��x���z1����1冚BIӱ�b�L9>>Pﶬ�/		IC}�;�Z�C.��]P;���'�[|����?�Pt���6w�^h�7Y��4��J��@aP?iE�42���f������94�����"C$s̫����5�P�=��õ�T^e�c�6�s�IBd���:멃H�(��ݶ��\m�#,Ec[��f��|;">�f��haUO��<e:ؤ�A��n�٭��D�����jV��<ƹ�p~Tj�oI>���d#�xЇA[`/T� �vTS ͜>\=un��=�{e�L��n�}�ؿ��fd,�?���^�% �t���t����R��>�@��Zu��a�=�>�||��~�~ݹ%�Q=�������kk �ޞq����G��\� ]4Jq���>~�f� m����1�e>q���4.���$�%A�/;���-�(9�+Y"�F���Wv��ǿ����T��T�v���'��!��Q����ʨ=��EU��a:��aYg�)l�� |A��~�晓�c��SUEE*��P�hn�#%m�_��+�H�`"��ӬPĽjW�)��݃q����iA�x�%JF�g�
?16.�z�
�W*��_`AD�97�f�fte�5��nq+��4��>��{־8Ϊ�cs��;x� �(a�*+��LC�����(��L�Mx(CCG�05�Ǯkl�w�p^+s�� b��ydhbb �|iee%j798D4u���<N�\���ڔ�Z�^N	g	"y��2��V�$�8:2���/G�;\?�r������䍐���J]�\��JKPDS�=H���ttb�����+����A���H��V�RQ��V��32x�ϷD)��i�X\��������	���t��:���q����4�,33�7#9��F�j��>B�e�g�&��[lj�3?77��xϾ�扣,�_��4X���

D�+4�j�IH�h�#Ӳk�;Ah�!���e}PD4��
'�����y�"�GD$��K�^�bOG��J�����%���9p|�8Ey�4|]�j�c����b���[3,��K���z�������ߔ��M�{�����3����~�)��gc��隙��C��n����-� ;��:�;_��t�{�'���X����Yɶ��|�Mgg�ys�8EH=kh%N&��>��]��Z�$OG��ȧo߾��6-p�)����哖�� F����~Ձ���F��x����,������}u�6����ҫL�r���@`��0񸆍���K@�����v�2�r
`��ǈKHX�-���uu!������Y��<�@Nb���I�.y�ß4���1I��¡q8�ؔ���@ZP#f�t��d�ț����T*F�W��~ffƈ�ɪ�����R��"�'��E�I0KKY�C`�94��3�OA#
�ң
<T_z����F󬭭G���FFF�4������ai�gb] [?����ly���8���|���D��b�n����\�ڐ,�a�����{6��WU�&>F6�QlƧ�A��Z�S����J�rq�IF`i��h���������}�ͩ �vA��A3 h419`YX���Ң�x�%i�ezJ�Y{ُ�Gv��u�u��q���4�}�MMM��u״C?}'jp�E���68m�LzON�OH���F VUU���N����r�΅WO�d\h����$.���\12<&�L2�|�x��9�ү��ik�
iȻ�R��������~��O�������8��k���ݸ:l�fAf�V��@w<M#�ZF���$$ܰ���MM�Zu��6F��Wd�Ӓ�z��LmN�������l�hs�Y�ǫ�LO����ұ����]��c�+W��ɷ��%�=����E�:,�,V���?1��n�UoH���y�з8����O�������R0k%!!qe�����A�ḻl`@���
b$rҡ�IG��bvu\TT��~�/uuu����ڻ'��h0!�~��aJ/`r�Xz?u�fJi��F�it�̇���`��z��z�����z���Y+�q'�f����$]@�(J��V����@{�������S��[}Ǵ�֦˲9M�ą������h���M�:##C��Q�8D�g�v!c4�b��(��S��������'�Y�W�G�L4kj:禧�)s���p�l?��gI�'c /����Bh��lR�D�� >���*jjBI}>�Ze��,r�[3@f��A^�L	����]hf.q�{����걖#�6L6��LY}�|�PW��.rB�k�-	r�\Xe�~�嘀S�)�0E� k����-ӳ�����1ܸ��22ζg���t0���"V�㰇����'O� �&�Wy���nl8�L�>=p���ňµ�BE4� ~�H�ݭ������Ϛ�v&��m��}���N� �AE����3�>}cy��.��W n���r�/G�p��s������i�N���7^o��E0Q��M--w��+��$��}U1��Ū<�姃��7(�(nj�W�����h_���-	�~�*��lh��,����� Ɂh\��x���3QM�CKg@�31.��lL�v��Ӥk��NG�>1&%����>_i(�R0��D����c�l��E�S�%me&�㝌�{Xb��u
� '���ƙ/�7iL,�&�ھ���˅�m�s��M�)���9Ki�ugc�˛��I��v���O�#<����MXA�B���8�c`v��Z�2Ѓ�͏������ݛ�ݩ��Ȟښ��q�r��呋���]	_���X��?�/k���)3��(��:������K��(�W�]޴Z�=�š����/*��%~���4:ON�}5�:G��{�W=x��-��t���Js��R1E�bb�kIN��Ϊ��p��{��R��+���xn����t7+��)��:�9B��C�iA�ZN��Iթ��̙��#C�R�y�������ЩE`�ȍ�±�b���u��/|��e���o�W�Z�C)�;X0�J_�  5�� �Y`�~�3$4Tz������h��&K �x�of�UV�L;s�% 5r]�}hd��B=�]�n�"b��ě����^�2{\>XO�/�p�/?������U����m���LV�] MEG�7XfZ]$\i{h�'|~qq1��V�H\2k:;��*�R�E*��C����ݬ�L����$	�x���_I��$VT����Sʠ.�}��E׾�6�����=ˤ�b�D�`�=�5|/�+���1�L�I�[y��/��~��(9qqq�>��aVIN����q��gϞͭn��t-�8/9~��)�[X�_{?�;)��`�A���­@&R��7G���]D~�P1��d��c���j��xᝐ�d*4�3DQ�FCJ�y�H�Y�n��K���hB�'�Y�iB��V��Y�J��.=��ο�:�9���^��Z�Y���=��ֳ�=��{�+�ӢEV����v���5h�::o";���^->&�d N���(���i`9L��?$"�W1�궏a����e�p�2����cv���N�����A�d����eG sl۶m<�yB�m$%�RF�1~~���N��iݘ��^�N���6�6�����Qm�~� 3"U+KK}��Cɜ^�|�wl�2-���
��n�_sm5�+R}~?ȭ]a;M���խjo���fXW��D[A!�� L^����✚o��C��1�Twg�h)��F���x�cn�ea3��V�ͫ�@�VS�=W�1[�6�(%Zn"V_V/�K�򼛛>T�ϕO��+v��!������י�������Q]�n�|�6H�Fz������|R2�x���2�v�{&����ì��/[��˫ԥ�ye�W�F����Tl����/_�/fa9�A��ݗu��X�=���@�� /�`|L䤕+Vt�F�}�m2[t����П�����!Oӷ�^��T��[�04���-U d'�t��C]�Yx���tR��f�J�)YPc5��@rr �̲]k��������R�ng��{�3г���H���]g%+���S�{�u�j���˭k��]]���
�9h���Z��~�E����P��~����$~���w^$RW[��������Bo�Ϗ��Mǖ�^2[��D�����?��u(�ſ��233���}��-fƓg��O�ך��>�����k�j�|�{��}zTz� �s5�U��?,����W��N���ލo���{{V-	R�q,Z1��P�DD1��B�T�#��܍Lc��:���+<�r~Oˏ������'O8�
p�y�n�֛fK����Ր>ׂ饾}T~�< h�@���C�� }3O�)z&�q��А���t�2H��7c�x���~��x%~�b����YR2��G�o՗I�F�˺�B��S^��`W��y��y���䏐�t�SP55�L�v�.�1~�-2 ����5�e9�YR��J�*�|G��l�6�Ns@MX����Ǫ�Ĭ�J����t������t�LR}�uѳ[�����,���l�	��@1ǽ����J�>FEw%V>���GZz:��C�E��8 ~�-�4褗����ֶR�_��nT��h���UE w���]��C?�!v>�n�d�C�k����z��s[��1Qo�<�5��_�	(*.����1V�t���k��FD�����O%j�/�@�K4f|||T
A���6��/�Q�XQud�\������
���n����@��-�IH$�%8�!*�9�uq�?A�u��	4��ޅ�S�$C�.�_YI]��g��gQ�@�r��
�PV��{M5�Q0�1��!I7�NI�RɃ�6�<�x��Zvvv�/���}�C�����QTTԣӑ������^/�7V���T��*J�ض�O|f#b�Zy�X���Ǡ��l�-�uu�ϕ� U��1����lr|�%ϽG��*9�����p/��}x�T�����>���Xy�&�h���l]Pv�\��#/^SZ�@Y�~�+d���t��0ק�Ŭ�[�8B��f͚5�����1�9�w~������Į��a`�i�*�3>%*3��~��Ԃ��4��*�"�MM�C��#TK�S�k�轭n�����\��U��J�.�jP,�����h�։V�ǿW�k����sr������f�̋-^[�>8%���f���D�V���!��_�O+**Z�b1����>�Q��_����g���v�C�~CƊN�_!Xn�����Y��uTħ�R��6�{��,�11뇃< Ӈ�QBq�q�{������X�<=#A��錭��!��#6�t����]>Y�4���W8Q�^	Y�E7���}���h��4L�P5�O�$�Ƞ:�9G��h唋�%nnn0�D"q�3�a��q�l��~�ePYW�L�ʚZ��ѥ?'��Ǎ�	(��z�<���q��b��:!��W���s�b��~�&7-��OnߌMi,פ����p��aze�U�.��¡L�	M#��F����c\��3��4X̽�Ƶ�.����V��K_��ж��w��&��{Oʏ�ܸq�WH�`ҟBϏ��|�����/���R�Fs�)�����r�	k��N�x�.�ĖKL "�F..��6q:,��z8��v:�Q��j$u��W^VG���t�D�}}^���܉k "��j7�?���ac�n~kz$�Y a\��Ũ�N��M8���%}�"�<�Sh��{�)m=@�κ��)��ҥ�k<�C�^�*fG���jV�����-�9@�E����Hス���ǏAm����Pz���Jn���#A�۸iSJ��j�i�Mר�h�d��|���e333Ә)����l�t1wN�w"�a�b~�g�t��|����ml,���~�4�KxB�m�-�ߵ��$~���c?��������=��|T����J���b�}�>�C�9� YR�k�*H��
���g'#����աq�.$���W�x,�VRR2�i���]5���u�t"�ENm�V��4�����g��p�Ѧ�"���8�)Z�B��ӛ�>��?�.��f��:���:�O���)�Sh/���=�����|����1�
�A(Gs�����zgQ���^ul�,9�n�~�0�������B��Ç����l���4����*n1{��C w���g�
÷��]�v�*���*�~|�

"�km�N�u��=Ŝ��,t$*�������,s��kEa	��O�v�:+�$m��o�}���ѱ�{����;��]�Gw<W���C��mrIގ66��Y��=i��:�H0�P<:s��`��dS&��N��ڨ�?1q���;��4�B=[���˗c�8�0I�"���nڅdY��q����Έ'O6@�������]vko�e�R@�I���*(�7�Q\^o}&���.�����H�S�5��Y(�])�}5L�iP���]��#;�w�ccբ7�~�Dgg��M�D_�h����RHTsg@�|Z�WE	 �!�"P"��\�vM0*H����6�F�_�<�o$���E�P�qM,���
*��+����&)�+�W�Y��U�F.�l��P|���T�[�FG�!oٰ���*���XdMŁce�WXL�
��``FT�f����Z�%��X\Q�_�8�Y@�Dhҿ�;i�5�	����Í�w��RE}�$K�0���Ϸ��ٛ�::��>�YI%B|�=��ܶ��0��&�7S�C��Ϫ��D~Z��8�,~�,����ɡ��R�hNʽ�:Ff�s
E#1)��]NZ�fJ���f0-������Z�xr�ӧ
L^�C��qt\�s.$w���� s����,�p�m�{g>Pu��صV��eܒ����4%�q<�t���^��EU�gve�������l��-����q�YN||�5#��O�[[/�5��
����m�\3n��_Մ:
27�|�����H�6.V� ���Q��e��F�u���0`�6&����಍1I������j$R�=nq���nxt��Kv*�kjjR/t�6bvoF/}��B�x9""���/j���|���R�:@G|L�]T���V 4X���<�t��#E�OZ��}� [__��[�wS 1������Ȏ
H8�3�65���:uwPYt�����t�BtC��kb��3{$���b��W�f�s\�,���&'#�M?����h=��[r_gō��2=lܾ����ﴒΓyw�.7��x߳zs����<��O����ٹ��'�f���_k�2�z�ȓ���q_>�:}�כKm��ٍ�ο/�l+5K��� &M�A/�v�e��Z�}�B�!�~o��5�ͬ�=;���E�t	ޮ��6T�O6Bexb��8���WUt�W]�b�ϟ?��탿C3�&�!.�{r/�K7H�H6̻g�H��XTL��\�0�1�hYhX�lt՝���b0/��ab����mTӼNO$�6��;�o<lڴI�wɛ���֢>?��R�&�������g�����5݃#���~ű�zw��*憫Q�<�����U  ���M����7�GR��7䲠��5��+ ٸ���o�+V���%C~<���DhI۸b�`��4��ArG,���f?����e��A'.�uX�;�=S=�������~d�P81��60 �$��<^�a5W�<V�5wV�%���g�n����b�Թ�"��^���G%�:��vH�A��W�o�� �.4���͛��Մ"��+۶�7�jI�����s�>� ���녚�����$W�U0=��F������{��N7\�1KEo����Rv0�� 0�\��Ӫ*M%�Ƣ\Qā��y�~��'�7����B,����v.Xk����j���F+�$��4y���BM��C������hD}oT����Xxcd؜2������孅�����������d��u�'�0������w�SbEm6�#5Q�r��g$�\�$ �_��X(27��'�Ӷ�l��1)f�ak"�{� �[9Ւ(0	��&��-4���M�����8��$\�i!/�9��:8:��? -zخ����yy�����������{5�_�*Iz�4<5ԭi'�fҤ�zC� ̈́B� �s5�e��C�o�C&����?�oMp�/J��-�2�Yfә��y���u+�����ՎX4�E���k����u����q5�AېQ�ɬ���<��e�MB�x��5ˍ�L����QuJ+�����%�o�OV�r7�n�4_@hX{"+;��g.^^���{�J�宵����6��U�����o�h�;�p�%i�� |`��r���Lw�<!.Vko�ת|�l��7%���N\\�4S2����@ݠ�X�|��6 �<f�k��3�%=%l�NzOH�e̴���HMZ�M�7�d���o�k�:�y�ff��=�e[��M�M:%iL���'m����$3C!��j���ߔ�G��4/����LP*&��#[�L[�|�� �u�U�;��{	B�0U?�iQ!��o�%�v�!�I#���C��=��O1������z999d ��V#�:�>I4�s^�о#a��Gž�<�Q�jo�#�B�D���ߎC\�m�x-tE�����"�����F��l��5ݑa��9�sG�V!e���헃�
[!����'HȅN���H����&���ڮ�v���P��TI=W��ۜ����$0���2���O��O��	���Aw��Z��m��Wq��s�F����*�!
���OW)	9gut�NR)�N4�ƊŞ�DpHXX�]��B��,�Ѵ��g̢�R'�$z�]d�z��qZ7��ll��1�������6��_� �p;v������t�fټf���>� I�9� ��Zvc��NـK��m�cŤ���=B�V,��-�'����߿���F߿Q��p3z�����|�351�hDI���ېEYXXl�]�J>�
>H௩L޽Y,e�����o�����ϛ�jo� �>�^��F�m���ݖ���h1X�䇢��4���2.��yr�ѴHک�|!�V�K�EFFV��<�tjj����WΏ��UyB�m�v//��h�������{'�"?��^�fS&靘��h�u���8�X�����ޓ����P��b�E�	;�~��� ����t��
to}	B���ӏW������_e>��G���A|m?�;��al�R��OK^��#1�~A��e����4_�$�='AX`�K3�$x�b�\��#q��3��=t ��
�������$�
�&ל��;t6�x��$t�%��ˣ{�Sp�h���>���% �?(s-�ԽbJ�L��q6\
�[/���*���H���*�hs<w�T�2�ߦ���e�"�����h�֢
��Z߹������/�t#;�˙��9��!���4�c=���if��}���c=}}E!�Z� ZH��mn��!Q��[��OQU�3w>$.���2s��XrTV� ���zo$��p%Y w�@��� �:�����f��=1118�g���i�/�il�T����D�n-m �>�N9��X�B2��ja[��"L�����%�J���O��\�����D䱁'`��Ā���/�{�b��v(?A�N#=:��h�ק-����қ���~��A���r�g��2%o��ܹ}e���tw	@��$H��s):���X��N��HKKS�Xв"�Z���*��I΁YP){����c7�y�c��D�����pby�ZrM!��=��� ߈Y���+�����F��Yc������2����@��������6/^���[����0�����9]\\^ggo�k�4�	&PUU��B��\7>���H�e�O!?<`�z��P��@h8=�.�lQ_�eCI:   �>��3�?p�^��v���雒r�7�O����`}���#@��\~~�S;#��橲���=(�!��8��
�%�w���{���S���$�w���;��;� @��O �u���ޮ��E���%� ������w]�zn���$'��#�h�]�Ҕڜ~�w�~�.@R<9���#P�Ԡj 4�yidd�U����Ք��j`��>A��[��AF�#j�!��C8L���*p%栍�a����w]�	� $F7�E����<�����Z(�`�U�fA��I�cp	���g;`�ɗ9r�|D�_/]�͜���H��RQGJDM:p/7�E�L���ӎ�v���Q�Ǖ(#��_�^F��|4V���C��y~�GHL���������;��]�=:���� �ֲ`�J�t�و�q��iH�M͏0f��"�7��E@�i�����aB(ף[��F�ggg�NIiSw�H~D�@��#w���'~3KE�p���X��#*@TK!%�5���!�T^F_f@��@&������,�ѯś�?�#D
�Ի
�84n6�#�IW���yHYzTy�+��
�Κ 2ˀg�JJ����D��u���@���r��\cJ��=߅�|SLR6�K�::���k�M�2�3��m��Ex��,u>H��@����@ ����T+��E�(f��t�������@�0׀oxX]�[-�V}���
K�6 ��+Qso�����E�Y���������fS�����U
i D�p��I~l.P�>�:V��\����t�[G�#��lZ�.̈́8�>����F�H7�8�$%M� ^������q�v�q��֓t�*I��*�<#@֐������n�K���Hˍ^�O�k ��W�R�fl�X&:��'������ad�]Uѯ32��_P�L6�ŷ�VVň����V�֜P,�eKǥQ��P�
ڛ��kH�sD I)\ʗ�L� ���n���S��߹[��n ��y|p22Ǘ�ߺit�u�7%K&:��\E�[vVn��R� ^ �|��ƿ���C��==�WzE�W!넄�>��1�V:���p��U:e
��O�i$ҿ���Ħ�êw��}�l-T���1�5f�K
�N1��zR�u��$==-]��d@=2�XI�!<<�f�./C��!���q�\�&�i�l6�������5��7�t��������_U�������\� $�E�<�]���"�<������t�廬d!�B��Uϡ��=(_Ƀ��^�'B�)��ucTkƯ�zݿ�.Giv0�Y	�--��`��F<�u`@Ŏ��p�F��^��BAY/L�y5J�|��-�x@���۵(�itH�c��Y+DPd�`F��Q�����q$�ҽ�%�c�h�&77���l$�)3�@��<���mX�=�	��sXpɐ�(��q�&����ۣbmpl��Dt�LdY�4Ru������:��)H���B���$���S 3��_(��Ӄ@/���$�ƅ�}�������MdQ2uuu�zrss��W>UA��V��'��s��ZL��_�ta�#�𽍖"����� ӏ���;{���Т_Z�z����L�i��������z�p�D{�ʻ�A��*Fx�/i[:i@��PՋX@�ԺLaj�f�A���ڌM��5� y����kz��~1vv�҈�f�R9����Li���+}j{�zbں5d�U��U~� P*d��VB���<$S��sj�|���r?@3���^����Ѹ��*:�����oL�h4��Ż�v����s\[O�U�"�u/��mP����/?�[(�$Z�����mT}�&�`%�T��e%��k0��Ç/XX����./�<$��$�M�':�P�zMl.m�M�F�В]˦PP*�
!�|/6cK����9Y��Z���'�6�'
�H�Kx6�~�ƿ>B5V�
�,�S��N\��zz��b��S�NA��������m��R,dK��h݉�D����3�\'�*�̱�q�y�[�Ys1�Q�A�(��8�C�jM۶��`oOK�t�re���c�]=��/�ӈ��6����c���9[jB����������Q��Zooo��,� ���'���(�Y�N�\1�Q�>�}�a�aE����C�Pa`1����X�r@5����Pg����m�C�9|Q4
���NCCw��!p��O�|뺶��MuU����V��]s�E�B�օPf�����WiƝ*�p�9�P�c����Pۻw/���Θ�������:G'*�iR��' �_�H ��L=�y��ә~
���z�ȏG�c�˰���2Ʉ�X�����󮀇 Ę��y��5��=$$� �����d-5QT�t;d���64����/��W@EĬ�e�M�6�'��9D�� �4Z�ԛ>�Ґ��ⶒW� �9��}����T@O�}R�����҅[����PG�S�w5��:��
��@��yANW�(��sp2����_��Z�	���4��
Ҏ�԰���;��37o��տ|�r�$��iG�n>0�}/@��$q�3	����Y�b~��Ŵ@��.���s���(��z��2��(��םṞ즡O�t/;�z���ʌ��}��95ONN����%�g�i��xH���$��t�4�����F_w����+��ď�y���OG&u����{�v��#[lA�`��QH�NÝ*��a�vV%Kq�Y��i�S��Y0�����pat *�rDq�66*l!�?�so�
�E&*x��;��èbho33=�?M��VA��ϠSȼy�" N��::��$5�Ԏ�L��hAC!aax��������
-�))�z��������VQ' 2���3�)�.���n��}Tcע/�@U���)��"�>h��0��w�m��l��}l��'�X��U����DQ@׀�燺��~f�� ͷA|E��u^�Իz�\�A9�@{ie!���^�9g!�F��-���N��V���m�����Pe�/נ?�EݧŪ $�
�h��o��Ѧ	�}[[�6-GA1e�Ж�7`����%�y�oDA4�J�܏J~��֡r�w��`�eAw�n�U��c�aO7��<H3Rh+
���$:�y�R? &HۈŹ�[���%��o��������C��h�җ��1��#	&z��h=L$-=�D���h&���Uu���9�!��բ
| |BϢ����������	�DM$C��qdn �3�M������+ShfP9i(J�l)������:����V�� ����𑲵��E2��xI���"�%�=��=��
��h��F��NII� ?��R~d�ٷ��[�r�Κ-��o[A���wݻ6l|���F�'1 �C5Z�S�6���NJ(Ix���px��+�6 %��_�~@�D��\"*���p�P�#�DA�~��̙3q����� �$�����Bݺ��V���`K ��� v� 7!�@?��}��IE���9#}�w��&d��Dx���@�/�w�}Z}�s�4l��!g�d���
=�C����γ�o�:m=�w>��}���`] \Q�z�"�� �@��
)�x�PA��-.ix�[�e�7�vȂ��s�� �����f���W���D����^DU[2-Oח��P�N�u���ٰ53�Dr���9h��6�_oq�ҽ
�/��;��Яs!G0x���iՒ�o������8��Z`��|XG`�[��+���Y�*v�*Fw�
,���m+����vvB����y�o~��l���$Rds!���
zO[-��W���&%GC" �!W���0Lu�F@��UY@��G��s����RT݃� �A� `A+ kNHN����`5��C`F[:���蘪	���`zE}�2y�������ޤ�K��������ab�A�Z�]ꍾ:ea��;-+k�4
|�m]�ȥ/R\�jq�2d����U�o�
�,T�� �DD�w��Ǡ0)�l�i�s��R	aL��i �/GNf��Y���hi���M~ŕ�U]�#��s�=����^[����P})PG|||���е�%���4A���谿���A/L��ҧ{n��� [��V���V2�oiu`c�@�[�%L�DFtA��\ 3h��H����}�>���~������6�mk�~�<�=�P��}���y���>�6���V�E��[�[9^ۥ|�l��X�~��haa!:������`���v5�b���`�ԃ� �4_-4�2���YX��W�Ջ����b@�M��!��T0`h*�c����㗟�[O��� ��7\���y;1O���X��TU}CCïz��e7?"ɒ�6(	`A��]�/}�xA���p����t5�p�r�>{l2�EŅ���̒t��/��M�h5��m���[����
w��/<��%,��7ȩ��&���=�F�y��������!ˬ½rBd_؇{Va�u܅&�5���fw��3kW"+�|L�:Eu$�Θ�>�3?�Q�Og))Qѱ�~��������͔���O�d����*������M{W�reZX �Μ�9τ����#�y3��M�,�#ˬɜlҦա%����S�h5,�:K���%�����深s�2�3|�h�V����c�(X}����%[Q zG4|M:sz(�;#7���A�8�h�8�]��K���,)�%CP;�1_��F\�8�^�uN�i`U�����!�Jg�:�Ƒ,C$��c$��^Dr5F�
H�. �Ia ��Eǥu0L\g�5��L��%xg���Z�L�4\����wFNM7�z6����K �
��;ܕ w
8��Owb�]
������0�>l���3�[��F���̓r=p�r��I�Ϛe��^��;�L���⦻���`��܋{R=	5p�r?� �I`�6��|�@=xX�ql�z�l��5�����Hr�Sn��-f��'�?�`�Ӡ�r�jue��?���A�Mw����,YƦ������VC�m0�P��П��p���:xă��<�'��I-�V�E��`����$�Q5B̳��k�����5)\P@�z�Y(���@�M'(�{�a̐��&�P#;��@O5��5�.V�F��Ƚ;-Y2��!l�<o�� ���&``���P��}Lj�,6�G7��;��)�}����ܛ�]?�3� ~�0�S��A��NO2�f� ^�d	�Q��1��la܂��:5�Ђ�p�B�Q����Hg;X�#(�I�,�U^"�ryբE_ާ�~yY~������	a�ˍ�'D��ě���n�7���^��bG�����%�7�~1�f�}�x����{��4/�bhc�'�lw�x�����<6݉��>�0�U��Ln#�}м [�aඃ�+>b�k6�d�~�m��}��,X����]�E���Q�o�Q���|�:v�(�K=�gZS��x��Jg.���0�\.���a��;��<Rs�9�`s�	�+�0F�B�� ږ>��C�%����дݡ����]�G��ׁ���8���@��9�3q���v)�tȶ���������J		=0OP�X+ a��9}�h����A�L��=A���ى�<�Q챫e�d�Ŏ8�_Q�I�Q.VL���jN_�7�=��+0�1�1��0#r �y`%6;s���6�[���+�n(ja%�b���0� ��-Xo?PhK��3��XC��8���P."�c*��jw �|�qr0=g��<��D���9Z^�q�8�1�uI�  ɂ� M{� .��b\�(�ԖJl6���<L{=�E�� �3B̯8����A[ڠ���V�A�F�Pg���A�0�!Ѝ��y��`�o�F����EY@:�X<�A*���C��zй�GN�1ȡ��=��������64��M�]n�`����uє7�O���d0�1x<z�P�I!xyV��z��<+-���j��G���!~@n+�ۍ�J��7���6z� <&�=�=���[�<�#��t.m*hT\[�=�6Nw���2kAL(�H�2��[��f�"��K�{Xg��,��)�A+`�3�rK.�� 3L���<��1���$�G�5�&*����a�%
3ʑ0иBἇ�\�t�� ���'���=��@�w�F1�-��߽��y9D���}�fl�ϐ���V��F&�̂�l�R.�}������Л#O�4�ڽ��]柈��-ւ��h�y��	���롣7p��!x,�ėNK;���z���Ή�)����߀��7���o����d�|��,������o�����?Tyß�m�$��q�M7�����W�v�(���(��%�mp���Zv%����.����)��<����1�R�25.����w���x�,�[������w$�R��@X%�����~�O^��v�����*���_ծ�1���#��9���F���,�o��l,Y�x���nof�Ϳ��:���������՛y����d!p�la��"�LK�:�I��v�\SS3���o:{��#:�rqq�`�s��U��\����w�ȴ�`k��+&ѻd��;��`N���І���C��&�ᶌE�mĕ�\W^�m̑'z�Z,�;z����&����f�u�3�8^��4�V�naU7����Q�*e@�1�
/PAGq)�-�w;,Y΁D�p��Jg�]���HB�}��gqcK�NgN��2|;<��eǵi��8g���4���ma�mÿ�o����2$.'����G�a
�Іی?z�ؠ���NÌq��|u��_7 ����m�9���^���#�����q���pM�ΞH����t��vVc�@�hÝ"��m��w:��NK�Nk����V#MK�[�vǷ�:��9������fh�yP~��ݲ�8ۑ%|]�Sja�q��Ƴ������#}a�7�3��mE�V�ZZ$U⒣��n罠��Pb���P �X/���FÃ!G�}�AA�����xP�]�{0�A��G�8	�S�Ծݚ%w< ����H<��=��u�ʊ����ߒ%ȟ�ݲ7�r9��P9T��n��Oa�5�!�ȴ�
.��~\Hp+L�6�nq�G��6�U�� �5@�G#XA&��0"����x���&���cp,���~���ha��Ex� �p���J�����v`j>�
��aj��=(^D�8FG5A��q<m7�m� ���Q$��ë��r���fl�0ƅ ����	�@n�	�����6�{���XW��~8�͒e	Lc�6�9���K���/��w��1�P"���k`���Jc�KnN��cx:� � ��Q__o����]ϴ`��v���?Y�$���q`�3fc-���i`w <�a
{ (�<�Jm���A��_ ,���n�%�e�EϘ��Ā�� �g츶�І�ۂk�!.߇��6D����6"zH�*�6D�w��:=����:��6f�m��D�������w������^_?�Ӕ��ǂ�ҟ0+7箯��y��E��������(�F�1�^� 2; 2��d���5�hǨ��D,�n��q�ȭ���]n����[,YZ$G4a�J"��Vk�� 1�� (�bFM�F�:�?`Ѓ��..lv���`dn�Hel����Գs0�	J=y�/=��a=n�`(�l#N���"�K�vূ�ԭ��у�@����"賥����v=�6(�C����{9@�W��a<A�@�ژ>3�e��(k�G��|sB�������2�B��`S� (9C1�W��NDp5Fp��>�wb���gG]]]C`>�!�%���b�3�][oς�bzр��J�`��w�L����T�
q��U^�D���Qah+��]�U��GU��]L2@O���6;�:���M~�; ��,Y�f����<"��Wɵ�}455���ߴn�q�EG��)�X6fa������bbډ(?��e��چ��xR���� z)y�$P`���*������	j�A��Sy9 ��0����R�|����� �P����c��)*6"h`��I��bn5����*�
� #ڸŚ�q��gv���-���P�ȳX�j|�k[�� s=;���$�`y&�z:,f+���0��5g��C뮑n�����c����%����|J��Rn�W��S�qmm�Xk]��̞fB�ۉ�����؟����F���c8}���|�Q��׌'�e�u���E�r���i�K<�$�Ý"�l���g:��%䌗|��Sd���c���D7C"����_$t�2��z�J�?}dE>�������Є�O2�����2���_���+�ꔈu���?+<
V���4�㿎��u��(ϑ�2��&�F��n5ޚ(�}}�ʢ��ݷ���V���\�S�^�����	��U]e՛(&f�O�}~v�Nv�Ԕ�?v�:^`m��v;d�jSM��#K���G'&���KM�.}�Y�<6�wf=�;@��j3o��?�N2��W�B��蠣�YV����c���7�A������p72�ѡΧU�5P5�ᨤ�&Y�ώ�d�mQg'5��Cՠ�i$��rO��믧����u�	h�E�'��1t�4�fK�R�k�{�>��A{���n�߄PR��$���I�T�W_=/�g�q`�{w�E>�LmB�"Rܙ�?��dN��q�ĭ#S[&������yǑ���\{��ә�C1��_�Y��/̮��aN=���d���=,&�!�a��"$�
�VX�ߜ"ߟҠ�����0q��lE�������h���T
��B�"�������B��_83h�DPVN�?�<�I�[��ş���*9C��Tiq�*T�|�����R�
U�lg`x�ƈX���t�r����x���wP�T�7v��A�aC�c#"����j�_�:TX&��hμs�g�Sf��w@�X#Z�/��ԟ��Z�P�i�y*E�"��k���4L5B���Kz�%�uӷw�7��v�t�,s9��WLE�7)ͺyvq����J�.?=���oi�xs���_?prk��k|��G}��a�
/+�C�ŚV��IDC��wޢk�2��ag�{��?Q1ȑ�����ԩ���mV�Hځ����>:S���'JL���3p�}P�O�?��zvh��l��=��V�Q-([G�a�\�^-ꬦ���u\i�@���-q*�z�2�T�Z����n@S�M�ۂg3��-)uFa�I؍Q��#���@3�pJ՞ZjW�����d�ԭ,���(��4�"�.�(ƻG�Ѷ%��c���,�!�!�9u&k�d�S�'�*�2�R��s/���zn"����Zo�|�d�5;4f���"���db�fMigف��$ܧ���k�f��>�x�?-)����I�y)b�N^���ՠb�㿨��ء��rxF��}*P\�雓�*�^v
��k9CU�.ػ�.�k���1pC�\x��v�eӡ�R��88#$)G(,q�Z$�����z�V�7L(��.���6���&n4�n]3���'�숓9�5rr�oRs(v������X��@���8ůT�%��o&>�S�0��R;�z�!�1�t���ܤ�
U\�a�m'��IԎ8Ǘ�����bQ��L&:��L�RT��_��F^�"n��ݺ��{a����xn�Ȝ�_���V%�N���U(�Dq�հJ������B�k��$��fe$��3x�����cмǌD��m4��Rg��UrS洄s��W�x���]V�$�H��տ�,Խ��&;�j�L¤���J������I�(���g�m�#F�|*�)�)��"��t���T��x�֦u�J�12��<�A�]��<�ϣ`�ie�'��W!�Lt~X���r���[TZ�ckB�ǉ��q�8#��Ó��s��?Qct䘼���JgS4F�8��w��eD��ΉC?�[iB�[tU�M�&>��^�넦Nn�w�7ڀ�o.�k��{{L��I���Pqd*ى�E�HjV��	�7����K,���E�k	�yo�L�mr/�-���Z_�jo�1Ev4�}�3fI���o����s�د��l�zpb7HW��E���eP�+r��z�)Vገ,�/6W�-)�������ɚ��Yo�?��4����(d@o��|�J@,{uo�h)�9�2@Q����ws�M�L�f�(�i3Pg�ӵ?ko��8�5bQȋ���Ϧҕ�Yv�r��HRS���ki�(���g�a  }��Ώ'Y�ޟ�|�ڞ?Ш{��M��X�$����K�����JN,O0P�yK<fok���lG�w���IW7��LH2[�Br�>���0Է?���SY�9�Q�r�VO�,����Z����씬����Ĕ���觢��r�r<�<.>:��T?��\Ú��H�g��2�zL\�yp}_1s�����Dt�K��3 	!5Z<��x���ZO���&��;���ニ:�}+u����1�T�<���/)+f�!"ݯrЎ�>�^��!2+͓�w&N:~DQ��T��)C��k��ҝr��UU�	��`B�wF�C�7yh�H�;�F�+�)�(�q�u�^�Xj��=�휾�L�0�����=����j���I>�xd4�,�)�lL|1����e�^��ߓ(u�����t��?��o�u���4��` ��3�&��b':x���'n
)^J쬾�('+#�]#�iYߦ�\��2:�� B�iTc���Zs��
/E���lg10��})u�a`D�Z�L!�E�J�O�� ���P����J��r�0���%ny�a8]�r���������0L�.+}\��?�c`�a%f��C�F.u�^� G����1Rg��r0v5ҍ	8�D|J��.�� �e`@:S��O�_�`@���������J�q��h�d�.�t�F߁=��=#:���Ga�?Ƶ�s���e��M�bYL����0!�<�R����d ��5�����\�\]�0��)�i��:ԟ�V�Iz���x�*��j���l��	�b`#=:V����g=��j�b��Q���<�~|��{��7�mUթv~ף�2�Ա�r������dz����NM�d@u�����b�Pg���ݓ\nka̾R8ձ(C��<���{��fٷK��� %����bf����K]�t�����qR�S�t2�g ��n�?��w�T�&yA��'m���F�~.��?�Ni�I���K��u�{oˀ��5iyq3:S?fy*f Q�3��U�u��������P�;��ș��Q�nC�72�zs������ݮ�e7��? ��>`W�-i\��:����6���!�7�m�����M��%���5�����c���Z�z��Aׯ��0&W��{���mP�7��]Kŗ�r2 ��rq�q���ͺn6O�̿i���#���l"#�?�g]x�e?���j!���z�VMjV���}#ī�|�^���K*��dEi���_�>8��4��:��`|w���	�K;V怳����(�W1��Qj���´��L�x���G��1"U�7��:�WԽ���ok��NPn&Z&5k4�;&��F�,܆����ɖ�3����rnvS5"Z�A�{�S^�m8�"Gef���.֐NsW2�f���?O\��;�_�`����
��4���F�)�,j�T��ԯ�}�3��a���Ru]���:N}�,�J�0\R�O��8w����1VZZZ.lN5gS��9���Z�=5<�;����;�đ�߇����E����Fø�/������d������s�����[�7���
�%zm��9�F�nJJ���I��T�ʹ�H��{`v��ѽ�\�NB�%�)�rr>2\}(�ִj�&��r5z�յ*��n��E`�O�Z��5N����@���~��ި���D)�)��oY7�j��rF������]��l�xy~�&Y�u�۝�3[�.A�ya��z��B����;[��X5�,�LS5����%5v�j�j�7�[�S�Sv�~ qb���늶�0�=������-w?�}N�p�	��M���2#�w�{��Ӝ݇�� �vt��Q��u��6jd���.��5i��R�6=�
���WIA��K9�YVBd�[�G)�#�(�{9W�UdI��fxh����'�U@b'C(u�R�r��S��,»7x��ʐ'~9:�fg��;����y$����:�oW(�(���yv9���Җ�Gmn/����6jZfZ�����	`�^r�F���̰#�U��v>v����L��Tg��a�MJ��+����I�f!⪄������i�I��bW�7k�c`I�E�C+�<�8�N���c�0^�p$��Ҭ:Ĭa:K��+�O�*3��u�Tza�d�3���)���AS�ī���?�t;Įo��e ;����k���mrl7����AkS���9�_��=71�$�Zu��ඳxBgH�a�)�u��R5�v���U=��[�f�FzY�s39��D|�:�\������X�º�:����q3J��x
�c0WY[{{Zyf���@�.^�¾Q/�O~�JcnW�Y��V�}O火K-�g)���,פ|Y�m�h�s�.�I?��Ԟa����"�2���s��F��w/.)�I��[��C�����B����Yi�m�@0W4�جW�A&�jC���Z�4�v��Û�1�<�D�ב_܆�Lx��*���5q���q���W#8���>_��ܾ�f,�]��G�c<Xte�i���:���5��%o2�X3�%��i*N\�-�%	Qk��;��z%o⽞ +QwD��OΏ'���#��Cuݜ�,�ň��*�JM��iۤ2;nQ��ab'�����x��db��#�������0/I�y��j�X%��q ��˰����K=8����`ͱ�׶�Ę��O����)��P��R��{�N�4�� ۵�ô���i��
�FŞ���"+�<��ˠ�o�o�T;s�N��63L�����J�먓����������"ý ��#o��j2���|L�C��`oo_�' zb�|·���
eѠ(f��n*ԡL�g��e�~2�U|b粰ӗ�9�2���/۫���8'yʱ1��\�꥕��v-ɻC���3_�EY)f�e����=����=����/h���+�Z��b��V�S7���K�gE@�!�"R@A�a	�X�֕Z[AP�%3!��HXԊ�7������|g��=��˽7s��O:j@!WN ��rDb�c�����Ȧ�0G��FI�ٮ��뮁\XBWxu.�L��,ۄm�߅�X�y3��W����_i�׻��ٸ��Y��v+�i;k��gd$O}T%�Ti;�7���]0Wft�O��w�J�5�����ѿUv���S&�nI"ҽӼx;�\����?ȱ�5k�d���C69��cUz���)l��&�f˜���ܥ^غ�*�N[����F�3��v�O�a�V9n�y��y����)����'�ކ�o���](C���m��{Yk{�禗w=ݕ8��n.����-{y����լ�Q��Ӕ����9G�\ࡴR)��G:�t|����e�&D�|�ѝ�;�Q�����.��
�5�YmVP��#�aa��d�֩Y��OSo�5d;�;V)5�cteI�n%���K���낌��C6��{AD;��$#c�_�ƒ~54��m��D���F��Z{��`�*��ȥjiGlXM�*�U����b{�"��	��fs��%������������k�g�+f���K���/���^�j�ϩE����K��s!>�/�/�j݉���k��8^��z�,���]WIxs�:B�q���dt�ő��Oޥ����'�����uȚ7��"��7|�KA�B2Ȗ78Gܲq{�$1C�Į~��8���v�B�u$=�I�<Ų�Q�w�,���gB�6��d�w#��_���re��<H����Ir(Rv+�Nw]}�x
9K�8�N��kJ��e�X}�F�r���*��D�֥x�؇Dڞ*A��s[[��9b�ӹax�б]�B�6-�ZR(3�a%��Ʃ���*{���j���6<��sE�A#���Un7_�k�6�U،����M��y?���|7�WP/�%��j��YD�9�=e�*�ڛ��;�mT�R��&y��F!��\���=O�(��>��q� G1A����Lk�������ӻ�kB���GtVd�_ݖj�B<��IcӇ�<yED�|º���TU���: {0�+�Я*OJ=x�DS��q����,x�m1:���K�<��@�3�x��6m�
9�.M�:7%y��[��-|�z��F���wW�e���%��C�k�ۻ�a���Gy��5�?8�hp)�3W��	��˜�k$��y{�|l9?��=�5�E�!��-ݎ��̎j}��@?���6ͪ]�����y�b2��!x��+/�$E�O�2�z2|Gz���r����{`���<��_1z�nq�/�ڎ�zU��}��������$[�/���������ks��Y�l���L������Ym���ԛĎ��o/�\hd�in��l9������G!b�#����&oN+(�إ#� ���\G���S������)���&�X��6S�LO!�X]�\I�����Ǥ�fo����eP���Й׏��рt>K����r6��t�ذYr?v���NӘ�@�<!�
5�'��+���p�N��^/��C���䌽<��R4� ���/ׁ��Q_�fɪ;y�分V��'�0,�����cǸi�Z�e�q�R]-2m�:�V �7O^ƍ�������<�\��=�K'��6[�_����������L�`t����f0�C��R�j�d��&E��c�o�D./��"=�hl�J��}U��(}��q�X8�xOc���!ٞ�>!M�J�h�N�(0G(�,$�񡬐�J�Z׍C�z|�Lѓ1�� �AY(�I�H�u�,q֥���B�X���m�bR/6�a��hm�k?��C��k�e��������^�7<t[?��uHorU��G�2�(s3D �3�rnpb�q:8ٖ��~wl}����5�c�
�����@�"KQ��P%�/O~��$Q/�w��<�y��tvǂ�=P�1��7Rk����z��Ɍ�"���C�ߙ����c�L5����=��O�*��̸oxH)/�
E���q��<�;���A^wQ^V0g��R&��@s(:{20G�xj��o�����=��yn��"��jO�a-X}12Y��L�K�����	1���c�j0#<Ʀ�LD�Į&�_*Ě;�zll������=%��iMf�a����w�s�6q�.�\��ԟ'���efG�H_�H�㖢x;�ĵlJ����J녲QG���i�4o�y���5Vg���O!_�Q�3V��T{fx� ?�ß���5�P��o�E��U)����-w W1��J�ŲQs˗9�uTU&u��<�(��z�`���7l��O���d��Z�xb*۴�{�{�)\��)�'[;���:�aB�Ui>�t��;�m��T�Ho�@g����)��$�x��ґ�e�u�=�&�����s�';r��y�AD'`�<d���EJB�;f=�H(��b�����K�$�"��D����vN/��XY����׋��8��C�f�˽%�#'�5lҨ'�m<���l�o2.�`e)SX/��R|͏���x�;�"Tẋ���0�N���֭���:��zFq ��]G���������w�Z�Ok|��W���an71������o�{Ug��
�}9"���!%��c��y��MᎵ���}�<�̍��(�sk�/�iAyv�Z�u��G*I�d�	��r�8W�.Pg�6`s�'�����:E�k�-"�r�[ ���s�����X9�S�����8�=��@:]�'�ZI(.�Pj����~����GDѮ��䑢A�h��4������z���F_�~��g�dsE�0G0x^�s)\�4����E��ѝ�����Uy�<Kv���y�D̋x;�!7[�^P�#���	k�4�d}��[݋�0�W޴��v��l}�\y�!�zA��x2�6��ƺ��%v�Q:[�=~� ���j�����T��y��5��~S�X�#t�����Vm�����K�&����������j7hp�+n��g�<�@�&���C�o	"�a���9Q�*�&+��,��8)��~`_k_m�Ȱ�΢�S��+�J���3� 2��J�m���h�}K�b]�Se`#�����Y˵��[�y�����?I
�`x�d��SQ3N�F�A��|S����ى����m�Zz�'<���BT��9ۿ�kc��;�*K�F�H,6!���/���9("��21������
o��E�~�f[1i�En�����aCD�!A��B�P�(�QTooRD��lT�^�}�
�|y{t�)�^E��8ޗ�f�#3LsĎD�Q�ݎl=u�1�l�ma��0MvY�$2�h]�O��a���Ǻ;�W�#��/�P�%{�����f��D�o��t_ $E�ě��"�$�o�W����Z#wҬ� i[ɞ�[�C�F�bu!C�/� "/FV_�)���P�9���y�l#�6�B��]g�p)����C�Z�\I[*�Eb=��}�6G��D�#ߚe���w5>��"2]��;��8��n$mɍ�ȩ]��Y���`���Yj�k� �ʔ�m�-E��Z�E0�ғ"�=[�?t��NA������a��U鈺�l�t_��k%�X@4A������Q �B����y�֓�Eg�U��go�e�}��-�����`��t��(s6ID�PF�ې�<�E�Q% %oDJ�C�_��j��Wp_��@��4y!�I<�/�<�k�-8�ҟH�m��Qfs�^�lYD��7L��@��]���rY%p����M$���1�m�P���T�^FX/�2�E��K�*ԗ����G|��v���Ԋu΢6�R��D��v(���G��R��FR0�9�%f]��5�.���靹���e��C���O��
z�㤠l�x��Z�Q�Ke�AE
W᎑��+.#-r}�Ґs�{n��g�~��ђ���%㇯����ﹿ�\}h�w"�J��Պw�SG��������Ӹv/��j�<\��k�!1�='t�����2ǻx�<<���?��p�O�E���t�(��M��?�&��Y�MG��&ǎڎ�!&	������G��È�-+-�o��.�o��ָ�YYI�]�Y7R��MN�:�_�1�tD���I��<��l���7��z�U���r�i�#j�l�buQ��*a� lo�5r�iQ���:�`��*��2�ʾ{�f�_�M	�݉}�LZ9-�m_���F��W����#��r��~{�N?�5�>8H7�7W}N�u�ٲ����N��ŁX�j��E�����+���c�:���� ��w����<_X%�����/��X�������= �v����z�,�� ���-��EB�����b;�D<R�Q"����]���x�҆�MT8&dT����&w���J�����D� �pn����%
��1@GR޼\����hG.���V`o�8n7� 
��7@NK&�ũ�3C�;����A�]��\ތ��k#�6��p�C��)=�)���
;ĳ��@�b�b�J��]��x��w�t��O�#�b���h�*܃��0�a��M9���,��?���Oq��zѦh��zn6،W��G�D;u�'�X�v���唂zD>��?!��m<��ؾ�m�~�Gj�[��W�R_�<���$b��s �NdJm�s�����e�"�ђ�D�U����[�Y� 6d+��a?� 
9O)=���&�U˚�lݎ�uHhd�?���"��Ȓ��9~*�=�8�͑�&�����H	�ž�B�V�]��S���s�Q�[����2^�٣]�k�19}r�����:r(e�^�W3@��Yӌ�L��Gz���T7P���5x���[,�`U%��*�As�u.[�v�z�˗-��:�Z}*�$cq�i��o{����SK���T}�I�ۦ��C�T޸1�� D�l�U���n��*&�������S�ۢ*����7������h��W�����)���HJ��i�5
}pT-���e3ƶ��I6���kp��
�[���؍���JuTY�O���	�[�>^�n�@sZ�����?O9�$�]/cZ;b�<]h�l��!d4@��{�����2~چy��8�����nha��YI_�c���Rh)�|r��ܐ����#���R���$�G���`W�v�y��eH,��ڲe�u遃H���6�'�0���5�J��!�8C�.��
��lC�9�0�	�}-��d#�Eٚ
:�x��(�~���S�ҌH�^q��Ą���p��c�����@��*֢�_GM�6���K���W"M�B	_I�İ��
u����*4��
v���PPXg�H�L�j/#g�s�Z���wD��|}1�AK,F+�#�JjĢq�m��
�������m�OG �\��,��RЃ^
NƟfD�Wz��^x�z!�U��;���r~�=����t�qҎ\�������U���+m��v)RZ��f��@��_��L�.�[G�aǅ��8�E��xV�"�V��U�$�"ϼv���p��!�_�q��x'#��E����\f'�_y�Opp�v!Z�GF����\T��[��v��O�v,�M]��zq��7��]�S���x�o2��i5���~�]�v�,�q��=�\@���x��<_���N�A�����R����p߶Szj��U��]�\ND߻�O��˟�W$45�.\��]���~�Tg��$6��,'�G�I�r��L�c�ωA�9�:G�C� ���3M,�0ݩ5H�ޤ��U�w��uE��|��vz��P�<�o�c���Tl)�Q~�l���ކ{�K�P�A������̃G�v��U���Ux�i#�el�Y��RQ$�%n��x�3�<����Uu�Y���+\\��R�/�Q���@�K�{��zZA�o�ޮ��f��2 7�`T��U��0\;��
-$���TH���]0���4#��B���?� &Ըq��]Y� b�Ĉ=X@����{�
3�u��4<�5�d���U5��`O�F�,<,�kTCS2*�Yf��b{0&��M�^'��.�@dg�WŽ����I��u��3V���۪j���N%F6���iʟW&Y��#��ۛ���ɼ�G�%�$Fv/@��lG"����K�#�B�ݗX��&�n�\DT���|�^(���yQ�3��V3���PQu!x�?���f3�A�z�w�&Uڒf�aѣ�.�V����ƕ��r�{I�qj,��~(B���0�Ryܦ4!Ʃy=G"YUH�[uƉAo���*ũ�I<�T�_�rـ�[���]=�V��V�����#�Wo���ǽz,�+=y�]uI���4Y��ǹ��o�'�-�kqA�$S�s�u7���D��O�X�c�B���ϭs�ղ)M��~���QBl�OꟌE�fC���,�VzcF�^� T"��v 9G]�6�}@�gVD5��U�.�9}Ű�F�
Ծh.�;��r���u�8m(����z��Ge�|���\d�D��r�	gۣ6��Q�b���H�����"+k~_"�l��Ȗ�әTH�(�c]�������0���[�g�x`�k��)8\5��C�t��*����ߍZ���\T�N�#L��I�o"w 5��>�D��|mr�K�S�������-h"���(�>�i>�d1�!���]6r�+�
���c��l�J���t�B���OX%�!$k��s�?���=]v^��a�ݔ36���.tw� �DH�Q ��U����C uM1x&��
r�M�\K�yj��u�N�ٺ�*�HU�L����r�8Q���\���b�3�?�v]���2�^���Ħ֮�ф���I����ee��벳K�dP��B/�!?]��&o򅎒i1��!�":��-QfH�b�֘Dċ5��f�����ش���^�����k�"��3��T�d�����~��(�Niag��� ��V6F쪮<
o��ȡyaO��XD؀?�FfDv��SB}��nL��#���D�q>����Bn�l5e�¡�D�c�҈�0�Er� %�������+}���fL�[*ۦ�};�:1�EB{�#j�&��ʑv�w���g���x�׋rĭ6��]� ��uNG.Æ*}7A�����s��}�LX���$�£ŋ���}B+y�.-d��T~��F��:�e`;�mV-�a©�F�J$�[����uK����m'D�ݧ{�a̭ƥQ՛s�N;B�3��j����2>���1 �Ͻtq�|�X|w�㟛�xr�TY�������|%��P lC��.3)$����^��Nb~�<�=*id�i�nd��UeKx>ԹI�t�"ד�rh���M�Z�]U�����U0�p�/[U�a��~�*S�G��.A��.���K$�X�|gD����k�R�)�&O[|q�w�kb1�in�r<L&���8E��G4�VkJ�&�^c�����m#�2M�Ew
C�*��+ݕ\����D��]K榋$^-5M�1�=��#���a1Dҍo^�cX�-�Co�!j�s���规��Gx���lI����)k/S��� W��{�E�*��h��~Dlo:��(�"M��h�������
m�`�I��RE�b�UuP�o����0�i(6��#'��5d�I݀�s?��W{U� ,�VU�|@�*����+�]����S�,����r��\ :GŐ�x\�^C�$c��j����W*�6i4\��{�����|M~v�*�G6"�K��cYˤ�ċI~��k���rrE��)��i��|�ZB֘:#�"�H�zMӐd�=7]`�P��K���D3��SV���7�&��S6s�Z�KG��h+���|�w�����f)_�s������I�����&����<2����׺z����؁H�qC80;����rF��L(�݌�6��r�e��^�z>���w�J��9���
:��p���dFBt,d�1��1#��,��i�g��md=��n�.G�7�{*��_~n��ly��c�A�&��z�/z�q�ŉ���9C#��g8\�5m?^�Iq0JC:P�@�mg=�Ƞz�Y/�3(C���A���+S"Y(�%d,XT� ��@���m���@y�E�F@iTz-f��`P�l*�r,( ]`=���
f���[Y���_�px���۾��Ȗ���t�	�Y7�%p���_t|>ޡ�!q@b[ k6�E�i��}��X@�5yhdBgȊ��:�tt�����]��`lN���/�
$�@M��d���=���KGZ�[�tX*���~�ʑ2S멜��O"bA?1F��N0H�������L(�H`�,�L'�Y>�H�r��:z)��� ��9R�eS �2Ћ�P�N`�^�7�Z �Ӟ�`��Џ28��~�o����xM IsA�
���z@e�ס�^�@���FA�^���6J��X�!%���]����r[��7�!!$ƜaL6~n����4۱4�����.�jP�{u�w+L\���E�Xyy��Ɵ���WCUg�{%��Zx-�J+��ZBs�O8��.�i�����?�eLǧ%'�^��bT���1�y��mF�4���]pu���FX,�~d`[X��`�F�f�ʂ1�,�Øq��.�>�X�V�_�Lj��}irh��!��>9Q�S{D��1=&%)�,S:5�q�ʑ�	{�>��n�6 �,f�- +e�΂l��lBg���j�ME��/�ě� �8���H�T ��R0#)���p�Mt�Ft�7��m�IFtp�2�����8�-�����T|A��4ͽg|�e�:�B-�4����t<0��H��?���':V|kdv�?���J�t�q��`7c�:;듟���� �ۓF�s��a�ǣ�FR)���-�n��h22�ĸ��P�s�m;M������ �m|�E0'_u���;��\T<Lw�������`�DEL(��f^�c\m���+� ��Oǀ�Mz�Vu,C@�;O�p��M ���`r���
~+�$�-��Z:�Rn�k0��3:eB8P8w�NS�gƅs�н���J�]�LHt4I6.���ӝ�|���h(:��h-��e�J�ke�o�ŧ+��
ş��`�Q�vC��@rAрQ��5 ���v��g2�0�p�s�av*H���OK-���`�!��Kx�w_�孍��k8��-�5h�`�c����44�g$������-&3
�f ��e�{���k�����i3_f��з"�C�|8�����į4`+A��v,�8��3�b�q ��'�0Gf���eƁ�ǟ6�x�8��	ֶ`��_��-��>n_7j3t$ �m5F���r.���΂?~�5�j��O�r��q�QT�����Qmw��	& ����/��5�3!���#��	G�m��杦�F�ݗ@z��{��Go�K�L�H��K���ß�- I�	R�$cC^V�$Y���?rC������޽�d޸����po��?2�[����r����PK   �v�X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   �v�X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   �v�X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   �v�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �v�X/yR�c  ^  /   images/d2af519c-c065-45b5-bffd-6bf239de2b90.png^��PNG

   IHDR   d   P   �	��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l��gw��c};��ΈU��ф#H�4�� �U�R����HU�V�z� �rD4��F��\���І�p8�Rb0�41���X������lf{vv����>�g��f�����������*�8ˏY&�d�xY���/�m\�BQ�6��#���a< )���������������~��f���rݟ���M�s���Ȳ���x= �IaB�� Zl�ۗ��������p�I���zV��ˊ������۷��v��/����,���$1�#L[ 	����t�ҥK���_����Y@NN�;wn�RRR�_s�â�Ͳ�e�[,>�7�AI�5DĐ�ˢ����I�&��2�M��	b���j����͇��cg��3,����r�x@c�0!W�\�[vG�p8���/���#�)��Qr��>��3L�9�e�OX6�FN�^(�1G����:joooHKK���"����.ܻ�e1�wYv��(�S/��t����P�������;D\I�Y��;,+YvRT���h�p�Ȼ�������Ғ3x�`b����M	��*�?�4�@�!�R�?x;��������/4A>��E�Yǲ�4W�{��(�ۉ	2n�8:~��~XŁ�Q��UWW�C��������Y^e��
&c�MFyy9�]��� e޼yqՏ�#)S��kg%���㏗s�=m���Ɋ+����
?o.?g3s��qLA��À�"V�k_�n]\�8�OI	���a��ڵk�9+2d9�N�&�|ʔ)t���)��@��<�zۇd)R�)���d�x���F�O��dgg��W2�T[[K���b�-�b�O�>B`�[�{������p�}RC&�6�gXo{�!��
b6o�L'N�S�N�p�]�}���Ni1w-�u ��ѣ�\�������h�ر4|�p��ʢ�S�Ү]���=�R��`8�)1���㡊�
�Ng�QSSC^�W([|���)4!H�"�T��u��bK�)wYY� %�� ���w������1		qdCo�B�p��R���L�'O�dXq;x�~��i6l�p�S���t����DEU#�)���y�2��SK��י �`\o���bU��1���@q� �Sc�����̌���A�Pt�K���7n�nJ�S ��Յb��[dS��o��f�q�V�Q��2(���]l}�4Q_?F�~l��=�������F���u8�)ܛ����R�2-�W�^d���is�uD�NXCC��5e6�u�LG+=9t�;؅����j������)/�y}����D�?蠃��G��M�L{��P�/�f�Iv[����-���p��N+�n A�&��y+')A�ج]J_�p�-�c\	N
̘1��/_N�������e��	VBA.�qd�̙��~I)h�v% [�Jo_�25ys�R���ug;=��h�����=[(1\���TO-���������tQ/+��2���Y�q,��!���l�U�������dy��V�WLt9����'��IA�0`�Ha�]�d	m߾�������`�cdn/��M�0!|��W�
f$�G�|���B�����a�r��.QN���E��S�e�l�t�(��9?�f�n$���,��4�jNO��"t$-�����A
Z<�pa�c�ܹsE9b\Z=������D2n��Ѱ���RЪ�����\A{/L�*�B߻<>l!�*զ)��qd�����.�a�7wO��n�f�=�<����nR'F���@�$��R��"�����/:yP<�-V�.�0ta �3���j-]����nѢ�lXHt�bq�C5����
�B�c�X݋Z|Y�V�T�����3�x� @]){��$�]`�� ��E"CF�v���`�޹�yp[pu�`�)�6�:�.�f����.�d@y(3[Ay�禋Q'��]U_	i�aAqA��ߣ�=�v~83"�{�V�,��1	]�p9P0������"�Bl!dVp] ���*�!��9���6_F�֔��Q�^�}(<�Z(�X'\n8}M��(
�Ҭ�4��2a!p;��mA�1z��gg �
��X#�fʰZ�Y�xϛ���1	ٸq#Z��髊1&��D�(n1&V�n��L�����Q���ƾUg�I��Ç�Q0��p�BJ��;!2�����X �C�Dn��ʕ+A�ZZZ�$J���28�T�y�f�}�>~ժUaRt%n0��TX�c<^!�,�IQ�u�����%�@�#�MT� ˈ�E'����6�=��z��B0�٤�H�L�w����!��	h����A���'�ǃ�	��SIH$�	뉢����!	��A�9�SS̰x�bw�@�u�������8����.��$���Y�9s����e˖)2�Jʃ>�zNN�M��֬"yܬHH�oD�F(�E�`�A[˒��e@�1;(1	n�[E�#�$����4���0xXPP�̟?_]�z���z%)2�?�p�\J�\��G��`���eI��X ����;��Z�;�x!ř� eŊ����ۡ[�СC�"p��c�xԨQʢE��M�6��d�HpV*^�q�UB?7�|������*���4�u$?PLՑ����<v��1hXb�q�̙1�����o�6��i)=�f�4к�:����yx?oڂ�0�����{����z<�=�-2#\�F�H�{���z	�~l����gY���O��h�uf0c�����>eVl}>�d��K�,ccU��P?z��k�Neǉ'�<�	E2vt����Ԏ��[�n5�V��$!�!:
����$B�/	I!��=ѧJY�"m9^,�!	Ijk{y��?��Kښa/��.*bJ�$$EX�tӫ���XxlK�dXb����t30��fڲs�ӣ�ZX�f	o�MZ/^ZH�C���늟���w�ÂD��&��$����38�MXXC��XK{5bU��O�諟It'0�T�vMu0Ȫ X����/�~¿"��t;LQ��'+}ݠ|>5�4��e?�v�߰%���?|饗���nX��,"-��;8��,{YvKBR��_+��wi.��1b�|IH
�ي��������_=�3�A��,��|��Q�\IH7C�)��+W�~��XO�e&��4ik�1�=����nF�UX�h�ol#�k��W�he�g����-$`��0���RFZF��F�e-���PW�`�ΨQ�^����>Â5��(�|6*<,	I�m�ǌ�>��e�|������,��V����ǉ�H�B���z�����_��V�B�0�.�|�4��$|��9IH
�q!n|���k�}bj�UB���9�X��]g�0�����V	��=�Y��D"��Κ�7�,dYb�|����$)�d@wm�����0)O��)B��fA���u�u��l��"��`���N���x�]?�~���&�e�_w:�x�$$�|��#G�|�ԩSq������A8c    IEND�B`�PK   �v�X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   �v�X�'k�  �  /   images/e8452abc-1b33-4025-a556-b46ce3c60df1.png��PNG

   IHDR   d   &   2r>3   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��[	�U��j{���zI��t0i�D���H$��3g<zt	G��AFe���(*3"�":.�
!,*[�$d![�ٺ�I��o����ߪ��@:�%��Mn���������zo��{r:�P$�����Jv�W��!�6Uuį��뚃�I�Op~�/���$�v�a�Pw��6�>j/��n���G�6�Tt��}l�St��~�S�J8���'����ċcÊ��h:��<���c�$�	�4@��}WM-M;0��Ј(��n�D�:��朵$��x���D����!G��t?���k�~�����]r��4�4��5��&E�NxO��i��}��\<�a&�9B�o�؈Ӹ�>�3+��ry�]T���C�ُ�ˏ@J�ìkA�e��(�϶��Έhϵ��3!��ܹ�!U�Ba�]�p!M�͜�'�Po!�8�I��sm���}瘊K��de��`?Sk�����^����i��P�"���b���LD�	��0/��ٔ��LB��:~b��*4��t����9�ae��"�K)Lȸ��t�y�GE[�e�I�Nc�W~d�⿎L}�B䉯���\a�d��V���5lL��1P]8
&]h$~�]�,��D���Wqd���t�p����1��jS�_[!b�tϣ X��B���cR�Z`�<X����2Ix��<ԧ,B�$1g�x��qV�.^��H������'N��B>�X�Dm}Y�ܰ�w�G�'f�y��h�2�r9H�	��gM��[�K_�aȧ��R�	է�fT(H��4 �^�&��P�j(Z
REx6TG�9LL1�z�RqZz4��A��"���jנ�	�W��U.P��m�ϩ��% W���ʑC�,&�� ��n#�D�j�Y��r�n����{�}�,`�@�f��I�|#̴i-T3n\>��щ�΀E�i�w$��� fϞ�k�����'.f���2A��A���~F0�'oCJ���(�Ť����j�Ѯ���h�v2�A�tt7��ۢ5I�+��>���� l^�;mC���v
%Ocڇ�N�!=z%�1���DL�����S�v���(�l�EA*�&��{;��ͨ8�MN:1t��P
�;��D� �?C�Waeft�Ǖ4�E��cČx@#f88�ȣ�&���iHU�h?�O?�$�.\H�I��4�2\��p` �H9�~�s;��/����a����0SK�*�a}V�g�F��b����&b�Al���j���A���o���	�]���VPtG�_~Ӆ�k�m���Q��`�ԃ�R��k����ކl�h���|F�5�����=�8O7����G�M����.�@�������G��Ryt&Iw؄h$	��":�%�>�Ïko��h�Q�1��H]y;ꪪn���K�޽�q0��Uo�`�RF����V�H�J�O�IT���Q�OP���$��"�
�L�k)/۵�8��6�I`ŭ�G����q8w��;y�y�������0=��D^��C��/K.,��E���4�T	�����]�<u�.���!��XJ��������7L̲ϙ�2����/���3���Y���1�"�L���%?_؞S&`�'��z�ʛl����9q,�"�d|�T	ӟ��4>��@���z�ۻ�%��!�m�w�Hr��A���+��@:�����A|���&�g����_��IÞ���u�1�y]���e�#PN"!�Q=�?��*b��;���j��i��Sf�R���F���,�aS0l��q��ڎ")(ɒ).��֧���p�Dmď�����t�CUdl>�Ep����i��5k��U��/�sd0��cv}�����m��xlk~E�wT��!̌A;�����R�o�pѠ�|-�WJ�xӨƄ�$:���H��X ym�E�R@��"����k$�:s y����1��fƺ]�8�>&^k�ϒ�G�X+�j���}�\��1�9g�^�eTo�z�`��}fnH������[qo�u���7&p��,_�4!E!�@���-˂��0MS<�w��4���4#&�>g�ْL1��]d35W"G��5̫���v�k*���֭_�K�/G�$���(b�`��T^����ά��C�;C�R�׆��Л"�9�Ag&���B��d�������4MS!Z]�444�
݋��ATWWc�̙hmmEKK��$:::��da|r��Wa�Q(`�h��Z��[�$DolCb������"�Yd�.��PY7�v*++a��0�����Khj�~�k�-|{;��e1C2��!L�

�V�x�Ј#VD0��e�SIn���V���)��kjj�`��Fz��؈T*�={���`�����*��ӧOǆ#q����c�k����y�SEL�H]&�%�m�=C͋������'��ޡ!��ރ��[a�*q�3����%��U����i��r</���l�\�.�ڱ
�)*&�E�ߧɱ:b5��:�Ţ`��g���+W
	:t������/b���طo���3Y\gFB-Y��&���M�@��*�dڞ>pS8�HӸ��B���a�����+?F�#�@	�g��N? 
&���h�˒</�k�M�;�I�ò��Ff!6Oɴ�
�^�7n��ȑ#BE]v�eصkv�܉ٳgU�u�Vq��ö�L[&~%<�� �-%�7�I"��Y��
I��
RY��W![�`���~�0�n���/aْ%�����˪��W���"����'�"�����F����Q�|j���N��Z�C���ǠdNڊ0CX-����Lٿ��f�Ē��mmm�%����=y�5Va����TY *Ո�
�j?yTgTI9�.�>2��:��[!�Ůh9��9�%��S�e-�z3�;<�� ���ݨ�6�*�Y �J���͛�x<���.tww�w�Vx��ѯ������8�3|4�O`*���0� �xW'�ɡfV�D�qp ���]��KR���6m:ló��a��������J�A��]/���"�ߎm c6��1���3��[UU%ο��jkk�!����bH$B���L{Y\�Btb�b�؅̈����	l��p2��$��E��� ��]���[��d%2��E���Q[Uq�/�o.�UV��@-_0����w�<<Sh&�0���l?]ac�c�aJd�ذ�
c;�##W�=X���0q�3���H�H*~��p�]����ds"�ۆV��ae�b [Q:k!�W}�?܃�tF��H_rl9���L���{�xte݄w�F�xU'��J�H�H8n�$�P��]��e�a/�$�y��R�2
KP]��Ϲ��zT$��y����Z�.���B!�-"g��/=$vk������G���éK9!�(/�=OpM�-��:VaO���,I�>	/�\Ċ��w�Q�Q��R��Ҕt���έ�A.o_�("���_{����}��f�~UxY%o?Čס>�?�{�~Z/���q��[��!��ea�Y�k��7L�QJd[.ֻpsh7μy����E��f(}�1¦,$r%�0�"�sk�¸�����J�w���.���_}��H]/k��4��T׌�6��؏.+�K��g����'��#��c���y�`{ ?�R�_T��X$5ў�(�.��l�Ķ�j�^�C[_��T=�����5/\��������tF}Rz��^� ������G���<E���L6V�L�퓧������;}-^'f�j�Ϛ �����EBIlPu�d�He�����8�)�𲊤�T�!�����?q�w ���#b�4�}b?$������p�|Z�P����8ht������K�N�ca���$�r�֏���<�t��,bjysJ<#��k8r�LT�,�h���y�}���Q,oCJ�_>4a{G�n [Qj�;�V�A�{�&�
U#���Zɡ\�����ק�e��gޫ�]C#�a�E���ӝi䟸��xj��` U<=b�;��7��[����f��:-���D�������8���i�i������.���7�v�rkx'��y�	xp�e=7	/��H}��I�v#u���҈؆��_T�lV�8���b/�S��i�dJ�ѕB`�;E|���t�b�e�q|Au�b�w0��f�3T��e$��׬���c΋#�s�nO������%�І^����\�d{!��Mqa�_h��u����"�4U�9�B)ً��F\r�%�'��
��kXa�&0�OQ]Hu�H.�=�c�əʹ�*���O���"����u����1(�%�"ͺ�3!�&�� ��V�~�Ex]i[��i.�[_���ދ�+V`��,�C��s0w��7�r�8O.2QC�	��/k��/�,sl���-�.X��Mq3�
�K�HNID�?�^>8(��_U����3�\9H�D��k��{�݇������-!�`(�_�����.��D�����J*k�)TV�038U���������,�����Nz۽�%�G���f�7�D��؉eq"��� ��N�6g{�,�Y#�!�Oo�}�ń�Kj��a��hy��]E#��}�uw�c�j[���_ �ę�4T�\�=uB�M8>l(5��%�&v�!�:�?�;�fy[Z�3�%�ENw�?�ݬ.80s�|���{~/G�!�a�����
Q��;q����#��A2�<�1Ln��a����,�8�p�p`J&���?��B�``�t]߲C'��v�Z�>D����ؒv�~X/ݏ�?܁���U������xO.�b��)J5ᛄ�§6>(����	o�q|�y�J��~��(8VKK���و�l,F3��S���.��	}��, ,i|�y��y��!�N�sv�z�"�N��&��k���l���a���z��#gaQ�ii� ���K�����6ࠀ�IZ!�#�l?����1��L�$�RQ��qR>>�ʛ#g�X���:1�[��&>�j��Hö�h~
2�e%&�e����P)��u�Øla���1#*�8gh&��
�wh}�P$Q��SDJݫ��d�"$	�f�CM�6(���K(�"�22�
��W@%��I�p#��C��E���-�?(#�Ȟ'ٌ����.t����)��B&<Z��:�'=~��Y��.�U�3�����!�P��yc�/�o/�]�����������I�nTV�q�G>5{�������pw׎HȤ�����>gP.V@|` ��r�	�L�0����2��~K�+R��"hOj5�U<X��dZ��O�L���:n�Bm��d�'��T�{��M铿I1�6[��`sp� f�DB�%��/#N�����a!1n!E��`��ջc=�q�}�����d��\���yMu�&�eq>kX-w2��b̟��HB�I����f��ؓ�ėV�G8R��FVF{�5�{r2"�#v�
�9��mT�H
�̔B��}ҲX�C��I�o��ICn�N8�.#k��;�2>�����6��Ǳ�`�!i˅� �]��f��q�](o��G����9�e��:Ё�S��*��b�|d��E���םX������)�؋)YT.<�<Mܻ�۽�M�W	�I�h�{�X�3��wƻ9#cS�]F|��w*�������������G������ß��go=<��c���79Gu�T�iT?�';T��G���Cf/�jJ�A&�	X������KD��'�o�
2�Iˆ��    IEND�B`�PK   �v�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �v�X	�I%�  �      jsons/user_defined.json��n���_E�Uh�9|���n������FQ��&*�
E���{%;�M�D�����F�Z3\߿f�/���2N���Ul~1�U���66����\������uCWӣ�}y�pjo��^�涆!޶�n>Ð�ٺ]��鯳��ɽ�Q��U�MK��r#��2"�EF����Q)�����c����M�l�Y=�_�N+Pn����W
#�(A���1U�2U,�+�ݲ��T��}�.��YW�5HUo�E۔0&��hmӾ�We�]��ۄU��iZH�q70V��0����3�8�\�+]7iz�6kX��u���U�_gé�\*��t�%,��Br��?��ln��fC�c
��l�4�6���#�Y����+S��9)W˅�|\/V��%;������;S�)�>��:��o�[�D�u���@m�x��'�K) 	��L���P=M��M[ރpO�j�6�Ö��e�Ad�����+�#܃m�����;�����v�\���K��^?�˦c�����b�j��o�Ml��bi��ZW/���O�*V��AX�{�ր��\.~��_�M=u���O�&��	<������7F�iP���	E��J�R�Q��%%� �yb�P

i*5�,XdC�(���O>z�^�:$-��j������ ��7�v�����`�@���d�y���6��J¥$�XH�s�~t?�}�1%��ݫ��Xy���Z°M	%�*d�6Hؖ��V_�ԫ&�j/�ɩ�Hd�a����6�$X������$�As�|��)rQ2�D
�r�������dU`�obU*��ɨ,�Nyd�qL�s����X��a1ySj뺽����}Jڛ��M�I�&�aqV;7�pf�b�-Oa�9ґ2D��vpV$����˴w6Y�y��v9�F�>j�I���vO��,�dJov�|��0�`\9R�icv��K��➾(�VDϸ����C���x��;�JV.����O�خ D�p��8���
 ��8j��E��� �"�����)0#���?�'w|�����]�	�QsA��@�CS�,<���y�C"/�=A�׶��br����rB���g࿯���v�n	�`H	u�r$��(z��pr�_=vcY'2Q�a3�����wY�� 
�`�p|��<B�@�X��Y��
)�#33�V�{�����<�}��F�
>�p�ڰ=5�*�*�8�unH!�ƺ� �	g�쉑�@�t�M@J��N`�)��K $T��P����Y�ӳ8��`c'p�����ˡ�cj�T�$G\i��*H] �ٗ}ބuYՓ��O�~W����ڦ^,�PNYp�c��)�aO��C�1���✎�<q41�tt�R*��9�>�rK�\�`�s8���Ѻ���OM!�ا�;:<l.gd�����ǋ���5�����
{sv������(���!M\��e�<�s�Q�"�9Ы�(�MΈʾ��ˢ��N�(�K���}Q:Jt������!�&ɗ�@3W�s��CE�U���E�H�q�?�y�>Pt\��E^�ϓ1xF���/���U��#eO�y���8��.$}���V���q�'dGq��"|�l:x,)���4-9V6�/t�i���&�:г�HU�W�3�q�1�*��g����2��Gl�ƨ�]��-6R5o�t�q�y��@�#U�t���%G���b�K�TŹ���K&�fy-���tB�i{w���>0��¿���e���+����˼q=�p���? PK
   �v�XiJʥ�  m�                   cirkitFile.jsonPK
   �v�X��(��8  �8  /               images/02932828-f6d4-4923-89fb-67d65ebd103a.pngPK
   �v�XR�\"# � /             7N  images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.pngPK
   �v�X� ���� 
� /             �q images/38cb4f51-bc72-4d24-b782-e5d855ce8001.pngPK
   �v�Xv��� f~ /             �( images/4d249bba-3190-4770-b321-fb8fc027a237.pngPK
   �v�X�1.:�  )  /             �0	 images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   �v�X?S��� 2� /             P	 images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   �v�X$�8�l  �  /             �' images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   �v�X$7h�!  �!  /             �E images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �v�X/yR�c  ^  /             �g images/d2af519c-c065-45b5-bffd-6bf239de2b90.pngPK
   �v�X�GDU7� �� /             �v images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   �v�X�'k�  �  /             -Z images/e8452abc-1b33-4025-a556-b46ce3c60df1.pngPK
   �v�XP��/�  ǽ  /             {q images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �v�X	�I%�  �                �# jsons/user_defined.jsonPK      �  �*   